/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: Multiplier_6_0_6_000

  Number system: Unsigned binary
  Multiplicand length: 7
  Multiplier length: 7
  Partial product generation: Simple PPG
  Partial product accumulation: Balanced delay tree
  Final stage addition: Brent-Kung adder
----------------------------------------------------------------------------*/

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_1(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_2(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_7(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_10(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_9(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_11(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_5(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_12(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_13_13(O);
  output [13:13] O;
  assign O[13] = 0;
endmodule

module GPGenerator(Go, Po, A, B);
  output Go;
  output Po;
  input A;
  input B;
  assign Go = A & B;
  assign Po = A ^ B;
endmodule

module CarryOperator(Go, Po, Gi1, Pi1, Gi2, Pi2);
  output Go;
  output Po;
  input Gi1;
  input Gi2;
  input Pi1;
  input Pi2;
  assign Go = Gi1 | ( Gi2 & Pi1 );
  assign Po = Pi1 & Pi2;
endmodule

module UBPriBKA_13_4(S, X, Y, Cin);
  output [14:4] S;
  input Cin;
  input [13:4] X;
  input [13:4] Y;
  wire [13:4] G0;
  wire [13:4] G1;
  wire [13:4] G2;
  wire [13:4] G3;
  wire [13:4] G4;
  wire [13:4] G5;
  wire [13:4] G6;
  wire [13:4] P0;
  wire [13:4] P1;
  wire [13:4] P2;
  wire [13:4] P3;
  wire [13:4] P4;
  wire [13:4] P5;
  wire [13:4] P6;
  assign P1[4] = P0[4];
  assign G1[4] = G0[4];
  assign P1[6] = P0[6];
  assign G1[6] = G0[6];
  assign P1[8] = P0[8];
  assign G1[8] = G0[8];
  assign P1[10] = P0[10];
  assign G1[10] = G0[10];
  assign P1[12] = P0[12];
  assign G1[12] = G0[12];
  assign P2[4] = P1[4];
  assign G2[4] = G1[4];
  assign P2[5] = P1[5];
  assign G2[5] = G1[5];
  assign P2[6] = P1[6];
  assign G2[6] = G1[6];
  assign P2[8] = P1[8];
  assign G2[8] = G1[8];
  assign P2[9] = P1[9];
  assign G2[9] = G1[9];
  assign P2[10] = P1[10];
  assign G2[10] = G1[10];
  assign P2[12] = P1[12];
  assign G2[12] = G1[12];
  assign P2[13] = P1[13];
  assign G2[13] = G1[13];
  assign P3[4] = P2[4];
  assign G3[4] = G2[4];
  assign P3[5] = P2[5];
  assign G3[5] = G2[5];
  assign P3[6] = P2[6];
  assign G3[6] = G2[6];
  assign P3[7] = P2[7];
  assign G3[7] = G2[7];
  assign P3[8] = P2[8];
  assign G3[8] = G2[8];
  assign P3[9] = P2[9];
  assign G3[9] = G2[9];
  assign P3[10] = P2[10];
  assign G3[10] = G2[10];
  assign P3[12] = P2[12];
  assign G3[12] = G2[12];
  assign P3[13] = P2[13];
  assign G3[13] = G2[13];
  assign P4[4] = P3[4];
  assign G4[4] = G3[4];
  assign P4[5] = P3[5];
  assign G4[5] = G3[5];
  assign P4[6] = P3[6];
  assign G4[6] = G3[6];
  assign P4[7] = P3[7];
  assign G4[7] = G3[7];
  assign P4[8] = P3[8];
  assign G4[8] = G3[8];
  assign P4[9] = P3[9];
  assign G4[9] = G3[9];
  assign P4[10] = P3[10];
  assign G4[10] = G3[10];
  assign P4[11] = P3[11];
  assign G4[11] = G3[11];
  assign P4[12] = P3[12];
  assign G4[12] = G3[12];
  assign P4[13] = P3[13];
  assign G4[13] = G3[13];
  assign P5[4] = P4[4];
  assign G5[4] = G4[4];
  assign P5[5] = P4[5];
  assign G5[5] = G4[5];
  assign P5[6] = P4[6];
  assign G5[6] = G4[6];
  assign P5[7] = P4[7];
  assign G5[7] = G4[7];
  assign P5[8] = P4[8];
  assign G5[8] = G4[8];
  assign P5[10] = P4[10];
  assign G5[10] = G4[10];
  assign P5[11] = P4[11];
  assign G5[11] = G4[11];
  assign P5[12] = P4[12];
  assign G5[12] = G4[12];
  assign P6[4] = P5[4];
  assign G6[4] = G5[4];
  assign P6[5] = P5[5];
  assign G6[5] = G5[5];
  assign P6[7] = P5[7];
  assign G6[7] = G5[7];
  assign P6[9] = P5[9];
  assign G6[9] = G5[9];
  assign P6[11] = P5[11];
  assign G6[11] = G5[11];
  assign P6[13] = P5[13];
  assign G6[13] = G5[13];
  assign S[4] = Cin ^ P0[4];
  assign S[5] = ( G6[4] | ( P6[4] & Cin ) ) ^ P0[5];
  assign S[6] = ( G6[5] | ( P6[5] & Cin ) ) ^ P0[6];
  assign S[7] = ( G6[6] | ( P6[6] & Cin ) ) ^ P0[7];
  assign S[8] = ( G6[7] | ( P6[7] & Cin ) ) ^ P0[8];
  assign S[9] = ( G6[8] | ( P6[8] & Cin ) ) ^ P0[9];
  assign S[10] = ( G6[9] | ( P6[9] & Cin ) ) ^ P0[10];
  assign S[11] = ( G6[10] | ( P6[10] & Cin ) ) ^ P0[11];
  assign S[12] = ( G6[11] | ( P6[11] & Cin ) ) ^ P0[12];
  assign S[13] = ( G6[12] | ( P6[12] & Cin ) ) ^ P0[13];
  assign S[14] = G6[13] | ( P6[13] & Cin );
  GPGenerator U0 (G0[4], P0[4], X[4], Y[4]);
  GPGenerator U1 (G0[5], P0[5], X[5], Y[5]);
  GPGenerator U2 (G0[6], P0[6], X[6], Y[6]);
  GPGenerator U3 (G0[7], P0[7], X[7], Y[7]);
  GPGenerator U4 (G0[8], P0[8], X[8], Y[8]);
  GPGenerator U5 (G0[9], P0[9], X[9], Y[9]);
  GPGenerator U6 (G0[10], P0[10], X[10], Y[10]);
  GPGenerator U7 (G0[11], P0[11], X[11], Y[11]);
  GPGenerator U8 (G0[12], P0[12], X[12], Y[12]);
  GPGenerator U9 (G0[13], P0[13], X[13], Y[13]);
  CarryOperator U10 (G1[5], P1[5], G0[5], P0[5], G0[4], P0[4]);
  CarryOperator U11 (G1[7], P1[7], G0[7], P0[7], G0[6], P0[6]);
  CarryOperator U12 (G1[9], P1[9], G0[9], P0[9], G0[8], P0[8]);
  CarryOperator U13 (G1[11], P1[11], G0[11], P0[11], G0[10], P0[10]);
  CarryOperator U14 (G1[13], P1[13], G0[13], P0[13], G0[12], P0[12]);
  CarryOperator U15 (G2[7], P2[7], G1[7], P1[7], G1[5], P1[5]);
  CarryOperator U16 (G2[11], P2[11], G1[11], P1[11], G1[9], P1[9]);
  CarryOperator U17 (G3[11], P3[11], G2[11], P2[11], G2[7], P2[7]);
  CarryOperator U18 (G5[9], P5[9], G4[9], P4[9], G4[7], P4[7]);
  CarryOperator U19 (G5[13], P5[13], G4[13], P4[13], G4[11], P4[11]);
  CarryOperator U20 (G6[6], P6[6], G5[6], P5[6], G5[5], P5[5]);
  CarryOperator U21 (G6[8], P6[8], G5[8], P5[8], G5[7], P5[7]);
  CarryOperator U22 (G6[10], P6[10], G5[10], P5[10], G5[9], P5[9]);
  CarryOperator U23 (G6[12], P6[12], G5[12], P5[12], G5[11], P5[11]);
endmodule

module UBZero_4_4(O);
  output [4:4] O;
  assign O[4] = 0;
endmodule

module Multiplier_6_0_6_000(P, IN1, IN2);
  output [13:0] P;
  input [6:0] IN1;
  input [6:0] IN2;
  wire [14:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  assign P[12] = W[12];
  assign P[13] = W[13];
  MultUB_STD_BLD_BK000 U0 (W, IN1, IN2);
endmodule

module BLDCON_8_2_8_0_11000 (S1, S2, IN0, IN1, IN2, IN3);
  output [12:3] S1;
  output [12:0] S2;
  input [8:2] IN0;
  input [8:0] IN1;
  input [11:5] IN2;
  input [11:3] IN3;
  wire [12:4] W1;
  wire [11:0] W2;
  CSA_8_0_11_5_11_3 U0 (W1, W2, IN1, IN2, IN3);
  CSA_12_4_11_0_8_2 U1 (S1, S2, W1, W2, IN0);
endmodule

module BLDTR_6_0_7_1_8_2000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6);
  output [13:4] S1;
  output [12:0] S2;
  input [6:0] PP0;
  input [7:1] PP1;
  input [8:2] PP2;
  input [9:3] PP3;
  input [10:4] PP4;
  input [11:5] PP5;
  input [12:6] PP6;
  wire [12:3] W0;
  wire [12:0] W1;
  BLDTR_6_0_7_1_8_2001 U0 (W0, W1, PP0, PP1, PP2, PP3, PP4, PP5);
  CSA_12_3_12_0_12_000 U1 (S1, S2, W0, W1, PP6);
endmodule

module BLDTR_6_0_7_1_8_2001 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5);
  output [12:3] S1;
  output [12:0] S2;
  input [6:0] PP0;
  input [7:1] PP1;
  input [8:2] PP2;
  input [9:3] PP3;
  input [10:4] PP4;
  input [11:5] PP5;
  wire [8:2] W0;
  wire [8:0] W1;
  wire [11:5] W2;
  wire [11:3] W3;
  UBARYACC_6_0_7_1_000 U0 (W0, W1, PP0, PP1, PP2);
  UBARYACC_9_3_10_4000 U1 (W2, W3, PP3, PP4, PP5);
  BLDCON_8_2_8_0_11000 U2 (S1, S2, W0, W1, W2, W3);
endmodule

module CSA_12_3_12_0_12_000 (C, S, X, Y, Z);
  output [13:4] C;
  output [12:0] S;
  input [12:3] X;
  input [12:0] Y;
  input [12:6] Z;
  UBCON_2_0 U0 (S[2:0], Y[2:0]);
  PureCSHA_5_3 U1 (C[6:4], S[5:3], X[5:3], Y[5:3]);
  PureCSA_12_6 U2 (C[13:7], S[12:6], Z[12:6], X[12:6], Y[12:6]);
endmodule

module CSA_12_4_11_0_8_2 (C, S, X, Y, Z);
  output [12:3] C;
  output [12:0] S;
  input [12:4] X;
  input [11:0] Y;
  input [8:2] Z;
  UBCON_1_0 U0 (S[1:0], Y[1:0]);
  PureCSHA_3_2 U1 (C[4:3], S[3:2], Z[3:2], Y[3:2]);
  PureCSA_8_4 U2 (C[9:5], S[8:4], X[8:4], Z[8:4], Y[8:4]);
  PureCSHA_11_9 U3 (C[12:10], S[11:9], X[11:9], Y[11:9]);
  UB1DCON_12 U4 (S[12], X[12]);
endmodule

module CSA_6_0_7_1_8_2 (C, S, X, Y, Z);
  output [8:2] C;
  output [8:0] S;
  input [6:0] X;
  input [7:1] Y;
  input [8:2] Z;
  UB1DCON_0 U0 (S[0], X[0]);
  UBHA_1 U1 (C[2], S[1], Y[1], X[1]);
  PureCSA_6_2 U2 (C[7:3], S[6:2], Z[6:2], Y[6:2], X[6:2]);
  UBHA_7 U3 (C[8], S[7], Z[7], Y[7]);
  UB1DCON_8 U4 (S[8], Z[8]);
endmodule

module CSA_8_0_11_5_11_3 (C, S, X, Y, Z);
  output [12:4] C;
  output [11:0] S;
  input [8:0] X;
  input [11:5] Y;
  input [11:3] Z;
  UBCON_2_0 U0 (S[2:0], X[2:0]);
  PureCSHA_4_3 U1 (C[5:4], S[4:3], Z[4:3], X[4:3]);
  PureCSA_8_5 U2 (C[9:6], S[8:5], Y[8:5], Z[8:5], X[8:5]);
  PureCSHA_11_9 U3 (C[12:10], S[11:9], Z[11:9], Y[11:9]);
endmodule

module CSA_9_3_10_4_11_5 (C, S, X, Y, Z);
  output [11:5] C;
  output [11:3] S;
  input [9:3] X;
  input [10:4] Y;
  input [11:5] Z;
  UB1DCON_3 U0 (S[3], X[3]);
  UBHA_4 U1 (C[5], S[4], Y[4], X[4]);
  PureCSA_9_5 U2 (C[10:6], S[9:5], Z[9:5], Y[9:5], X[9:5]);
  UBHA_10 U3 (C[11], S[10], Z[10], Y[10]);
  UB1DCON_11 U4 (S[11], Z[11]);
endmodule

module MultUB_STD_BLD_BK000 (P, IN1, IN2);
  output [14:0] P;
  input [6:0] IN1;
  input [6:0] IN2;
  wire [6:0] PP0;
  wire [7:1] PP1;
  wire [8:2] PP2;
  wire [9:3] PP3;
  wire [10:4] PP4;
  wire [11:5] PP5;
  wire [12:6] PP6;
  wire [13:4] S1;
  wire [12:0] S2;
  UBPPG_6_0_6_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, IN1, IN2);
  BLDTR_6_0_7_1_8_2000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6);
  UBBKA_13_4_12_0 U2 (P, S1, S2);
endmodule

module PureCSA_12_6 (C, S, X, Y, Z);
  output [13:7] C;
  output [12:6] S;
  input [12:6] X;
  input [12:6] Y;
  input [12:6] Z;
  UBFA_6 U0 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U1 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U2 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U3 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U4 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U5 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U6 (C[13], S[12], X[12], Y[12], Z[12]);
endmodule

module PureCSA_6_2 (C, S, X, Y, Z);
  output [7:3] C;
  output [6:2] S;
  input [6:2] X;
  input [6:2] Y;
  input [6:2] Z;
  UBFA_2 U0 (C[3], S[2], X[2], Y[2], Z[2]);
  UBFA_3 U1 (C[4], S[3], X[3], Y[3], Z[3]);
  UBFA_4 U2 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U3 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U4 (C[7], S[6], X[6], Y[6], Z[6]);
endmodule

module PureCSA_8_4 (C, S, X, Y, Z);
  output [9:5] C;
  output [8:4] S;
  input [8:4] X;
  input [8:4] Y;
  input [8:4] Z;
  UBFA_4 U0 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U1 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U2 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U3 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U4 (C[9], S[8], X[8], Y[8], Z[8]);
endmodule

module PureCSA_8_5 (C, S, X, Y, Z);
  output [9:6] C;
  output [8:5] S;
  input [8:5] X;
  input [8:5] Y;
  input [8:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U3 (C[9], S[8], X[8], Y[8], Z[8]);
endmodule

module PureCSA_9_5 (C, S, X, Y, Z);
  output [10:6] C;
  output [9:5] S;
  input [9:5] X;
  input [9:5] Y;
  input [9:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U3 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U4 (C[10], S[9], X[9], Y[9], Z[9]);
endmodule

module PureCSHA_11_9 (C, S, X, Y);
  output [12:10] C;
  output [11:9] S;
  input [11:9] X;
  input [11:9] Y;
  UBHA_9 U0 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U1 (C[11], S[10], X[10], Y[10]);
  UBHA_11 U2 (C[12], S[11], X[11], Y[11]);
endmodule

module PureCSHA_3_2 (C, S, X, Y);
  output [4:3] C;
  output [3:2] S;
  input [3:2] X;
  input [3:2] Y;
  UBHA_2 U0 (C[3], S[2], X[2], Y[2]);
  UBHA_3 U1 (C[4], S[3], X[3], Y[3]);
endmodule

module PureCSHA_4_3 (C, S, X, Y);
  output [5:4] C;
  output [4:3] S;
  input [4:3] X;
  input [4:3] Y;
  UBHA_3 U0 (C[4], S[3], X[3], Y[3]);
  UBHA_4 U1 (C[5], S[4], X[4], Y[4]);
endmodule

module PureCSHA_5_3 (C, S, X, Y);
  output [6:4] C;
  output [5:3] S;
  input [5:3] X;
  input [5:3] Y;
  UBHA_3 U0 (C[4], S[3], X[3], Y[3]);
  UBHA_4 U1 (C[5], S[4], X[4], Y[4]);
  UBHA_5 U2 (C[6], S[5], X[5], Y[5]);
endmodule

module UBARYACC_6_0_7_1_000 (S1, S2, PP0, PP1, PP2);
  output [8:2] S1;
  output [8:0] S2;
  input [6:0] PP0;
  input [7:1] PP1;
  input [8:2] PP2;
  CSA_6_0_7_1_8_2 U0 (S1, S2, PP0, PP1, PP2);
endmodule

module UBARYACC_9_3_10_4000 (S1, S2, PP0, PP1, PP2);
  output [11:5] S1;
  output [11:3] S2;
  input [9:3] PP0;
  input [10:4] PP1;
  input [11:5] PP2;
  CSA_9_3_10_4_11_5 U0 (S1, S2, PP0, PP1, PP2);
endmodule

module UBBKA_13_4_12_0 (S, X, Y);
  output [14:0] S;
  input [13:4] X;
  input [12:0] Y;
  wire [13:4] Z;
  UBExtender_12_4_1000 U0 (Z[13:4], Y[12:4]);
  UBPureBKA_13_4 U1 (S[14:4], X[13:4], Z[13:4]);
  UBCON_3_0 U2 (S[3:0], Y[3:0]);
endmodule

module UBCON_12_4 (O, I);
  output [12:4] O;
  input [12:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
  UB1DCON_11 U7 (O[11], I[11]);
  UB1DCON_12 U8 (O[12], I[12]);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBCON_3_0 (O, I);
  output [3:0] O;
  input [3:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
endmodule

module UBExtender_12_4_1000 (O, I);
  output [13:4] O;
  input [12:4] I;
  UBCON_12_4 U0 (O[12:4], I[12:4]);
  UBZero_13_13 U1 (O[13]);
endmodule

module UBPPG_6_0_6_0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, IN1, IN2);
  output [6:0] PP0;
  output [7:1] PP1;
  output [8:2] PP2;
  output [9:3] PP3;
  output [10:4] PP4;
  output [11:5] PP5;
  output [12:6] PP6;
  input [6:0] IN1;
  input [6:0] IN2;
  UBVPPG_6_0_0 U0 (PP0, IN1, IN2[0]);
  UBVPPG_6_0_1 U1 (PP1, IN1, IN2[1]);
  UBVPPG_6_0_2 U2 (PP2, IN1, IN2[2]);
  UBVPPG_6_0_3 U3 (PP3, IN1, IN2[3]);
  UBVPPG_6_0_4 U4 (PP4, IN1, IN2[4]);
  UBVPPG_6_0_5 U5 (PP5, IN1, IN2[5]);
  UBVPPG_6_0_6 U6 (PP6, IN1, IN2[6]);
endmodule

module UBPureBKA_13_4 (S, X, Y);
  output [14:4] S;
  input [13:4] X;
  input [13:4] Y;
  wire C;
  UBPriBKA_13_4 U0 (S, X, Y, C);
  UBZero_4_4 U1 (C);
endmodule

module UBVPPG_6_0_0 (O, IN1, IN2);
  output [6:0] O;
  input [6:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
  UB1BPPG_6_0 U6 (O[6], IN1[6], IN2);
endmodule

module UBVPPG_6_0_1 (O, IN1, IN2);
  output [7:1] O;
  input [6:0] IN1;
  input IN2;
  UB1BPPG_0_1 U0 (O[1], IN1[0], IN2);
  UB1BPPG_1_1 U1 (O[2], IN1[1], IN2);
  UB1BPPG_2_1 U2 (O[3], IN1[2], IN2);
  UB1BPPG_3_1 U3 (O[4], IN1[3], IN2);
  UB1BPPG_4_1 U4 (O[5], IN1[4], IN2);
  UB1BPPG_5_1 U5 (O[6], IN1[5], IN2);
  UB1BPPG_6_1 U6 (O[7], IN1[6], IN2);
endmodule

module UBVPPG_6_0_2 (O, IN1, IN2);
  output [8:2] O;
  input [6:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
  UB1BPPG_6_2 U6 (O[8], IN1[6], IN2);
endmodule

module UBVPPG_6_0_3 (O, IN1, IN2);
  output [9:3] O;
  input [6:0] IN1;
  input IN2;
  UB1BPPG_0_3 U0 (O[3], IN1[0], IN2);
  UB1BPPG_1_3 U1 (O[4], IN1[1], IN2);
  UB1BPPG_2_3 U2 (O[5], IN1[2], IN2);
  UB1BPPG_3_3 U3 (O[6], IN1[3], IN2);
  UB1BPPG_4_3 U4 (O[7], IN1[4], IN2);
  UB1BPPG_5_3 U5 (O[8], IN1[5], IN2);
  UB1BPPG_6_3 U6 (O[9], IN1[6], IN2);
endmodule

module UBVPPG_6_0_4 (O, IN1, IN2);
  output [10:4] O;
  input [6:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
  UB1BPPG_6_4 U6 (O[10], IN1[6], IN2);
endmodule

module UBVPPG_6_0_5 (O, IN1, IN2);
  output [11:5] O;
  input [6:0] IN1;
  input IN2;
  UB1BPPG_0_5 U0 (O[5], IN1[0], IN2);
  UB1BPPG_1_5 U1 (O[6], IN1[1], IN2);
  UB1BPPG_2_5 U2 (O[7], IN1[2], IN2);
  UB1BPPG_3_5 U3 (O[8], IN1[3], IN2);
  UB1BPPG_4_5 U4 (O[9], IN1[4], IN2);
  UB1BPPG_5_5 U5 (O[10], IN1[5], IN2);
  UB1BPPG_6_5 U6 (O[11], IN1[6], IN2);
endmodule

module UBVPPG_6_0_6 (O, IN1, IN2);
  output [12:6] O;
  input [6:0] IN1;
  input IN2;
  UB1BPPG_0_6 U0 (O[6], IN1[0], IN2);
  UB1BPPG_1_6 U1 (O[7], IN1[1], IN2);
  UB1BPPG_2_6 U2 (O[8], IN1[2], IN2);
  UB1BPPG_3_6 U3 (O[9], IN1[3], IN2);
  UB1BPPG_4_6 U4 (O[10], IN1[4], IN2);
  UB1BPPG_5_6 U5 (O[11], IN1[5], IN2);
  UB1BPPG_6_6 U6 (O[12], IN1[6], IN2);
endmodule

