/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: Multiplier_11_0_9000

  Number system: Unsigned binary
  Multiplicand length: 12
  Multiplier length: 10
  Partial product generation: Simple PPG
  Partial product accumulation: Dadda tree
  Final stage addition: Han-Carlson adder
----------------------------------------------------------------------------*/

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UBHA_9(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_12(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_6(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_7(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_8(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_12(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_13(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_14(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_15(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_5(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_16(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_17(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_18(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_19(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module GPGenerator(Go, Po, A, B);
  output Go;
  output Po;
  input A;
  input B;
  assign Go = A & B;
  assign Po = A ^ B;
endmodule

module CarryOperator(Go, Po, Gi1, Pi1, Gi2, Pi2);
  output Go;
  output Po;
  input Gi1;
  input Gi2;
  input Pi1;
  input Pi2;
  assign Go = Gi1 | ( Gi2 & Pi1 );
  assign Po = Pi1 & Pi2;
endmodule

module UBPriHCA_20_1(S, X, Y, Cin);
  output [21:1] S;
  input Cin;
  input [20:1] X;
  input [20:1] Y;
  wire [20:1] G0;
  wire [20:1] G1;
  wire [20:1] G2;
  wire [20:1] G3;
  wire [20:1] G4;
  wire [20:1] G5;
  wire [20:1] G6;
  wire [20:1] P0;
  wire [20:1] P1;
  wire [20:1] P2;
  wire [20:1] P3;
  wire [20:1] P4;
  wire [20:1] P5;
  wire [20:1] P6;
  assign P1[1] = P0[1];
  assign G1[1] = G0[1];
  assign P1[3] = P0[3];
  assign G1[3] = G0[3];
  assign P1[5] = P0[5];
  assign G1[5] = G0[5];
  assign P1[7] = P0[7];
  assign G1[7] = G0[7];
  assign P1[9] = P0[9];
  assign G1[9] = G0[9];
  assign P1[11] = P0[11];
  assign G1[11] = G0[11];
  assign P1[13] = P0[13];
  assign G1[13] = G0[13];
  assign P1[15] = P0[15];
  assign G1[15] = G0[15];
  assign P1[17] = P0[17];
  assign G1[17] = G0[17];
  assign P1[19] = P0[19];
  assign G1[19] = G0[19];
  assign P2[1] = P1[1];
  assign G2[1] = G1[1];
  assign P2[2] = P1[2];
  assign G2[2] = G1[2];
  assign P2[3] = P1[3];
  assign G2[3] = G1[3];
  assign P2[5] = P1[5];
  assign G2[5] = G1[5];
  assign P2[7] = P1[7];
  assign G2[7] = G1[7];
  assign P2[9] = P1[9];
  assign G2[9] = G1[9];
  assign P2[11] = P1[11];
  assign G2[11] = G1[11];
  assign P2[13] = P1[13];
  assign G2[13] = G1[13];
  assign P2[15] = P1[15];
  assign G2[15] = G1[15];
  assign P2[17] = P1[17];
  assign G2[17] = G1[17];
  assign P2[19] = P1[19];
  assign G2[19] = G1[19];
  assign P3[1] = P2[1];
  assign G3[1] = G2[1];
  assign P3[2] = P2[2];
  assign G3[2] = G2[2];
  assign P3[3] = P2[3];
  assign G3[3] = G2[3];
  assign P3[4] = P2[4];
  assign G3[4] = G2[4];
  assign P3[5] = P2[5];
  assign G3[5] = G2[5];
  assign P3[7] = P2[7];
  assign G3[7] = G2[7];
  assign P3[9] = P2[9];
  assign G3[9] = G2[9];
  assign P3[11] = P2[11];
  assign G3[11] = G2[11];
  assign P3[13] = P2[13];
  assign G3[13] = G2[13];
  assign P3[15] = P2[15];
  assign G3[15] = G2[15];
  assign P3[17] = P2[17];
  assign G3[17] = G2[17];
  assign P3[19] = P2[19];
  assign G3[19] = G2[19];
  assign P4[1] = P3[1];
  assign G4[1] = G3[1];
  assign P4[2] = P3[2];
  assign G4[2] = G3[2];
  assign P4[3] = P3[3];
  assign G4[3] = G3[3];
  assign P4[4] = P3[4];
  assign G4[4] = G3[4];
  assign P4[5] = P3[5];
  assign G4[5] = G3[5];
  assign P4[6] = P3[6];
  assign G4[6] = G3[6];
  assign P4[7] = P3[7];
  assign G4[7] = G3[7];
  assign P4[8] = P3[8];
  assign G4[8] = G3[8];
  assign P4[9] = P3[9];
  assign G4[9] = G3[9];
  assign P4[11] = P3[11];
  assign G4[11] = G3[11];
  assign P4[13] = P3[13];
  assign G4[13] = G3[13];
  assign P4[15] = P3[15];
  assign G4[15] = G3[15];
  assign P4[17] = P3[17];
  assign G4[17] = G3[17];
  assign P4[19] = P3[19];
  assign G4[19] = G3[19];
  assign P5[1] = P4[1];
  assign G5[1] = G4[1];
  assign P5[2] = P4[2];
  assign G5[2] = G4[2];
  assign P5[3] = P4[3];
  assign G5[3] = G4[3];
  assign P5[4] = P4[4];
  assign G5[4] = G4[4];
  assign P5[5] = P4[5];
  assign G5[5] = G4[5];
  assign P5[6] = P4[6];
  assign G5[6] = G4[6];
  assign P5[7] = P4[7];
  assign G5[7] = G4[7];
  assign P5[8] = P4[8];
  assign G5[8] = G4[8];
  assign P5[9] = P4[9];
  assign G5[9] = G4[9];
  assign P5[10] = P4[10];
  assign G5[10] = G4[10];
  assign P5[11] = P4[11];
  assign G5[11] = G4[11];
  assign P5[12] = P4[12];
  assign G5[12] = G4[12];
  assign P5[13] = P4[13];
  assign G5[13] = G4[13];
  assign P5[14] = P4[14];
  assign G5[14] = G4[14];
  assign P5[15] = P4[15];
  assign G5[15] = G4[15];
  assign P5[16] = P4[16];
  assign G5[16] = G4[16];
  assign P5[17] = P4[17];
  assign G5[17] = G4[17];
  assign P5[19] = P4[19];
  assign G5[19] = G4[19];
  assign P6[1] = P5[1];
  assign G6[1] = G5[1];
  assign P6[2] = P5[2];
  assign G6[2] = G5[2];
  assign P6[4] = P5[4];
  assign G6[4] = G5[4];
  assign P6[6] = P5[6];
  assign G6[6] = G5[6];
  assign P6[8] = P5[8];
  assign G6[8] = G5[8];
  assign P6[10] = P5[10];
  assign G6[10] = G5[10];
  assign P6[12] = P5[12];
  assign G6[12] = G5[12];
  assign P6[14] = P5[14];
  assign G6[14] = G5[14];
  assign P6[16] = P5[16];
  assign G6[16] = G5[16];
  assign P6[18] = P5[18];
  assign G6[18] = G5[18];
  assign P6[20] = P5[20];
  assign G6[20] = G5[20];
  assign S[1] = Cin ^ P0[1];
  assign S[2] = ( G6[1] | ( P6[1] & Cin ) ) ^ P0[2];
  assign S[3] = ( G6[2] | ( P6[2] & Cin ) ) ^ P0[3];
  assign S[4] = ( G6[3] | ( P6[3] & Cin ) ) ^ P0[4];
  assign S[5] = ( G6[4] | ( P6[4] & Cin ) ) ^ P0[5];
  assign S[6] = ( G6[5] | ( P6[5] & Cin ) ) ^ P0[6];
  assign S[7] = ( G6[6] | ( P6[6] & Cin ) ) ^ P0[7];
  assign S[8] = ( G6[7] | ( P6[7] & Cin ) ) ^ P0[8];
  assign S[9] = ( G6[8] | ( P6[8] & Cin ) ) ^ P0[9];
  assign S[10] = ( G6[9] | ( P6[9] & Cin ) ) ^ P0[10];
  assign S[11] = ( G6[10] | ( P6[10] & Cin ) ) ^ P0[11];
  assign S[12] = ( G6[11] | ( P6[11] & Cin ) ) ^ P0[12];
  assign S[13] = ( G6[12] | ( P6[12] & Cin ) ) ^ P0[13];
  assign S[14] = ( G6[13] | ( P6[13] & Cin ) ) ^ P0[14];
  assign S[15] = ( G6[14] | ( P6[14] & Cin ) ) ^ P0[15];
  assign S[16] = ( G6[15] | ( P6[15] & Cin ) ) ^ P0[16];
  assign S[17] = ( G6[16] | ( P6[16] & Cin ) ) ^ P0[17];
  assign S[18] = ( G6[17] | ( P6[17] & Cin ) ) ^ P0[18];
  assign S[19] = ( G6[18] | ( P6[18] & Cin ) ) ^ P0[19];
  assign S[20] = ( G6[19] | ( P6[19] & Cin ) ) ^ P0[20];
  assign S[21] = G6[20] | ( P6[20] & Cin );
  GPGenerator U0 (G0[1], P0[1], X[1], Y[1]);
  GPGenerator U1 (G0[2], P0[2], X[2], Y[2]);
  GPGenerator U2 (G0[3], P0[3], X[3], Y[3]);
  GPGenerator U3 (G0[4], P0[4], X[4], Y[4]);
  GPGenerator U4 (G0[5], P0[5], X[5], Y[5]);
  GPGenerator U5 (G0[6], P0[6], X[6], Y[6]);
  GPGenerator U6 (G0[7], P0[7], X[7], Y[7]);
  GPGenerator U7 (G0[8], P0[8], X[8], Y[8]);
  GPGenerator U8 (G0[9], P0[9], X[9], Y[9]);
  GPGenerator U9 (G0[10], P0[10], X[10], Y[10]);
  GPGenerator U10 (G0[11], P0[11], X[11], Y[11]);
  GPGenerator U11 (G0[12], P0[12], X[12], Y[12]);
  GPGenerator U12 (G0[13], P0[13], X[13], Y[13]);
  GPGenerator U13 (G0[14], P0[14], X[14], Y[14]);
  GPGenerator U14 (G0[15], P0[15], X[15], Y[15]);
  GPGenerator U15 (G0[16], P0[16], X[16], Y[16]);
  GPGenerator U16 (G0[17], P0[17], X[17], Y[17]);
  GPGenerator U17 (G0[18], P0[18], X[18], Y[18]);
  GPGenerator U18 (G0[19], P0[19], X[19], Y[19]);
  GPGenerator U19 (G0[20], P0[20], X[20], Y[20]);
  CarryOperator U20 (G1[2], P1[2], G0[2], P0[2], G0[1], P0[1]);
  CarryOperator U21 (G1[4], P1[4], G0[4], P0[4], G0[3], P0[3]);
  CarryOperator U22 (G1[6], P1[6], G0[6], P0[6], G0[5], P0[5]);
  CarryOperator U23 (G1[8], P1[8], G0[8], P0[8], G0[7], P0[7]);
  CarryOperator U24 (G1[10], P1[10], G0[10], P0[10], G0[9], P0[9]);
  CarryOperator U25 (G1[12], P1[12], G0[12], P0[12], G0[11], P0[11]);
  CarryOperator U26 (G1[14], P1[14], G0[14], P0[14], G0[13], P0[13]);
  CarryOperator U27 (G1[16], P1[16], G0[16], P0[16], G0[15], P0[15]);
  CarryOperator U28 (G1[18], P1[18], G0[18], P0[18], G0[17], P0[17]);
  CarryOperator U29 (G1[20], P1[20], G0[20], P0[20], G0[19], P0[19]);
  CarryOperator U30 (G2[4], P2[4], G1[4], P1[4], G1[2], P1[2]);
  CarryOperator U31 (G2[6], P2[6], G1[6], P1[6], G1[4], P1[4]);
  CarryOperator U32 (G2[8], P2[8], G1[8], P1[8], G1[6], P1[6]);
  CarryOperator U33 (G2[10], P2[10], G1[10], P1[10], G1[8], P1[8]);
  CarryOperator U34 (G2[12], P2[12], G1[12], P1[12], G1[10], P1[10]);
  CarryOperator U35 (G2[14], P2[14], G1[14], P1[14], G1[12], P1[12]);
  CarryOperator U36 (G2[16], P2[16], G1[16], P1[16], G1[14], P1[14]);
  CarryOperator U37 (G2[18], P2[18], G1[18], P1[18], G1[16], P1[16]);
  CarryOperator U38 (G2[20], P2[20], G1[20], P1[20], G1[18], P1[18]);
  CarryOperator U39 (G3[6], P3[6], G2[6], P2[6], G2[2], P2[2]);
  CarryOperator U40 (G3[8], P3[8], G2[8], P2[8], G2[4], P2[4]);
  CarryOperator U41 (G3[10], P3[10], G2[10], P2[10], G2[6], P2[6]);
  CarryOperator U42 (G3[12], P3[12], G2[12], P2[12], G2[8], P2[8]);
  CarryOperator U43 (G3[14], P3[14], G2[14], P2[14], G2[10], P2[10]);
  CarryOperator U44 (G3[16], P3[16], G2[16], P2[16], G2[12], P2[12]);
  CarryOperator U45 (G3[18], P3[18], G2[18], P2[18], G2[14], P2[14]);
  CarryOperator U46 (G3[20], P3[20], G2[20], P2[20], G2[16], P2[16]);
  CarryOperator U47 (G4[10], P4[10], G3[10], P3[10], G3[2], P3[2]);
  CarryOperator U48 (G4[12], P4[12], G3[12], P3[12], G3[4], P3[4]);
  CarryOperator U49 (G4[14], P4[14], G3[14], P3[14], G3[6], P3[6]);
  CarryOperator U50 (G4[16], P4[16], G3[16], P3[16], G3[8], P3[8]);
  CarryOperator U51 (G4[18], P4[18], G3[18], P3[18], G3[10], P3[10]);
  CarryOperator U52 (G4[20], P4[20], G3[20], P3[20], G3[12], P3[12]);
  CarryOperator U53 (G5[18], P5[18], G4[18], P4[18], G4[2], P4[2]);
  CarryOperator U54 (G5[20], P5[20], G4[20], P4[20], G4[4], P4[4]);
  CarryOperator U55 (G6[3], P6[3], G5[3], P5[3], G5[2], P5[2]);
  CarryOperator U56 (G6[5], P6[5], G5[5], P5[5], G5[4], P5[4]);
  CarryOperator U57 (G6[7], P6[7], G5[7], P5[7], G5[6], P5[6]);
  CarryOperator U58 (G6[9], P6[9], G5[9], P5[9], G5[8], P5[8]);
  CarryOperator U59 (G6[11], P6[11], G5[11], P5[11], G5[10], P5[10]);
  CarryOperator U60 (G6[13], P6[13], G5[13], P5[13], G5[12], P5[12]);
  CarryOperator U61 (G6[15], P6[15], G5[15], P5[15], G5[14], P5[14]);
  CarryOperator U62 (G6[17], P6[17], G5[17], P5[17], G5[16], P5[16]);
  CarryOperator U63 (G6[19], P6[19], G5[19], P5[19], G5[18], P5[18]);
endmodule

module UBZero_1_1(O);
  output [1:1] O;
  assign O[1] = 0;
endmodule

module Multiplier_11_0_9000(P, IN1, IN2);
  output [21:0] P;
  input [11:0] IN1;
  input [9:0] IN2;
  wire [21:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  assign P[12] = W[12];
  assign P[13] = W[13];
  assign P[14] = W[14];
  assign P[15] = W[15];
  assign P[16] = W[16];
  assign P[17] = W[17];
  assign P[18] = W[18];
  assign P[19] = W[19];
  assign P[20] = W[20];
  assign P[21] = W[21];
  MultUB_STD_DAD_HC000 U0 (W, IN1, IN2);
endmodule

module DADTR_11_0_12_1_1000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9);
  output [20:0] S1;
  output [20:1] S2;
  input [11:0] PP0;
  input [12:1] PP1;
  input [13:2] PP2;
  input [14:3] PP3;
  input [15:4] PP4;
  input [16:5] PP5;
  input [17:6] PP6;
  input [18:7] PP7;
  input [19:8] PP8;
  input [20:9] PP9;
  wire [20:0] W0;
  wire [19:1] W1;
  wire [18:2] W2;
  wire [17:3] W3;
  wire [16:4] W4;
  wire [15:5] W5;
  wire [14:6] W6;
  wire [13:7] W7;
  wire [13:8] W8;
  UBHA_9 U0 (W7[10], W8[9], PP0[9], PP1[9]);
  UBFA_10 U1 (W7[11], W8[10], PP0[10], PP1[10], PP2[10]);
  UBFA_11 U2 (W7[12], W8[11], PP0[11], PP1[11], PP2[11]);
  UBHA_12 U3 (W8[13], W8[12], PP1[12], PP2[12]);
  UBCON_8_0 U4 (W0[8:0], PP0[8:0]);
  UB1DCON_9 U5 (W0[9], PP2[9]);
  UBCON_12_10 U6 (W0[12:10], PP3[12:10]);
  UB1DCON_13 U7 (W0[13], PP2[13]);
  UB1DCON_14 U8 (W0[14], PP3[14]);
  UB1DCON_15 U9 (W0[15], PP4[15]);
  UB1DCON_16 U10 (W0[16], PP5[16]);
  UB1DCON_17 U11 (W0[17], PP6[17]);
  UB1DCON_18 U12 (W0[18], PP7[18]);
  UB1DCON_19 U13 (W0[19], PP8[19]);
  UB1DCON_20 U14 (W0[20], PP9[20]);
  UBCON_8_1 U15 (W1[8:1], PP1[8:1]);
  UB1DCON_9 U16 (W1[9], PP3[9]);
  UBCON_12_10 U17 (W1[12:10], PP4[12:10]);
  UB1DCON_13 U18 (W1[13], PP3[13]);
  UB1DCON_14 U19 (W1[14], PP4[14]);
  UB1DCON_15 U20 (W1[15], PP5[15]);
  UB1DCON_16 U21 (W1[16], PP6[16]);
  UB1DCON_17 U22 (W1[17], PP7[17]);
  UB1DCON_18 U23 (W1[18], PP8[18]);
  UB1DCON_19 U24 (W1[19], PP9[19]);
  UBCON_8_2 U25 (W2[8:2], PP2[8:2]);
  UB1DCON_9 U26 (W2[9], PP4[9]);
  UBCON_12_10 U27 (W2[12:10], PP5[12:10]);
  UB1DCON_13 U28 (W2[13], PP4[13]);
  UB1DCON_14 U29 (W2[14], PP5[14]);
  UB1DCON_15 U30 (W2[15], PP6[15]);
  UB1DCON_16 U31 (W2[16], PP7[16]);
  UB1DCON_17 U32 (W2[17], PP8[17]);
  UB1DCON_18 U33 (W2[18], PP9[18]);
  UBCON_8_3 U34 (W3[8:3], PP3[8:3]);
  UB1DCON_9 U35 (W3[9], PP5[9]);
  UBCON_12_10 U36 (W3[12:10], PP6[12:10]);
  UB1DCON_13 U37 (W3[13], PP5[13]);
  UB1DCON_14 U38 (W3[14], PP6[14]);
  UB1DCON_15 U39 (W3[15], PP7[15]);
  UB1DCON_16 U40 (W3[16], PP8[16]);
  UB1DCON_17 U41 (W3[17], PP9[17]);
  UBCON_8_4 U42 (W4[8:4], PP4[8:4]);
  UB1DCON_9 U43 (W4[9], PP6[9]);
  UBCON_12_10 U44 (W4[12:10], PP7[12:10]);
  UB1DCON_13 U45 (W4[13], PP6[13]);
  UB1DCON_14 U46 (W4[14], PP7[14]);
  UB1DCON_15 U47 (W4[15], PP8[15]);
  UB1DCON_16 U48 (W4[16], PP9[16]);
  UBCON_8_5 U49 (W5[8:5], PP5[8:5]);
  UB1DCON_9 U50 (W5[9], PP7[9]);
  UBCON_12_10 U51 (W5[12:10], PP8[12:10]);
  UB1DCON_13 U52 (W5[13], PP7[13]);
  UB1DCON_14 U53 (W5[14], PP8[14]);
  UB1DCON_15 U54 (W5[15], PP9[15]);
  UBCON_8_6 U55 (W6[8:6], PP6[8:6]);
  UB1DCON_9 U56 (W6[9], PP8[9]);
  UBCON_12_10 U57 (W6[12:10], PP9[12:10]);
  UB1DCON_13 U58 (W6[13], PP8[13]);
  UB1DCON_14 U59 (W6[14], PP9[14]);
  UBCON_8_7 U60 (W7[8:7], PP7[8:7]);
  UB1DCON_9 U61 (W7[9], PP9[9]);
  UB1DCON_13 U62 (W7[13], PP9[13]);
  UB1DCON_8 U63 (W8[8], PP8[8]);
  DADTR_20_0_19_1_1000 U64 (S1, S2, W0, W1, W2, W3, W4, W5, W6, W7, W8);
endmodule

module DADTR_20_0_19_1_1000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8);
  output [20:0] S1;
  output [20:1] S2;
  input [20:0] PP0;
  input [19:1] PP1;
  input [18:2] PP2;
  input [17:3] PP3;
  input [16:4] PP4;
  input [15:5] PP5;
  input [14:6] PP6;
  input [13:7] PP7;
  input [13:8] PP8;
  wire [20:0] W0;
  wire [19:1] W1;
  wire [18:2] W2;
  wire [17:3] W3;
  wire [16:4] W4;
  wire [16:5] W5;
  UBHA_6 U0 (W3[7], W5[6], PP0[6], PP1[6]);
  UBFA_7 U1 (W1[8], W4[7], PP0[7], PP1[7], PP2[7]);
  UBHA_7 U2 (W2[8], W5[7], PP3[7], PP4[7]);
  UBFA_8 U3 (W0[9], W3[8], PP0[8], PP1[8], PP2[8]);
  UBFA_8 U4 (W1[9], W4[8], PP3[8], PP4[8], PP5[8]);
  UBHA_8 U5 (W2[9], W5[8], PP6[8], PP7[8]);
  UBFA_9 U6 (W0[10], W3[9], PP0[9], PP1[9], PP2[9]);
  UBFA_9 U7 (W1[10], W4[9], PP3[9], PP4[9], PP5[9]);
  UBFA_9 U8 (W2[10], W5[9], PP6[9], PP7[9], PP8[9]);
  UBFA_10 U9 (W0[11], W3[10], PP0[10], PP1[10], PP2[10]);
  UBFA_10 U10 (W1[11], W4[10], PP3[10], PP4[10], PP5[10]);
  UBFA_10 U11 (W2[11], W5[10], PP6[10], PP7[10], PP8[10]);
  UBFA_11 U12 (W0[12], W3[11], PP0[11], PP1[11], PP2[11]);
  UBFA_11 U13 (W1[12], W4[11], PP3[11], PP4[11], PP5[11]);
  UBFA_11 U14 (W2[12], W5[11], PP6[11], PP7[11], PP8[11]);
  UBFA_12 U15 (W0[13], W3[12], PP0[12], PP1[12], PP2[12]);
  UBFA_12 U16 (W1[13], W4[12], PP3[12], PP4[12], PP5[12]);
  UBFA_12 U17 (W2[13], W5[12], PP6[12], PP7[12], PP8[12]);
  UBFA_13 U18 (W1[14], W3[13], PP0[13], PP1[13], PP2[13]);
  UBFA_13 U19 (W2[14], W4[13], PP3[13], PP4[13], PP5[13]);
  UBFA_13 U20 (W3[14], W5[13], PP6[13], PP7[13], PP8[13]);
  UBFA_14 U21 (W3[15], W4[14], PP0[14], PP1[14], PP2[14]);
  UBFA_14 U22 (W4[15], W5[14], PP3[14], PP4[14], PP5[14]);
  UBFA_15 U23 (W5[16], W5[15], PP0[15], PP1[15], PP2[15]);
  UBCON_5_0 U24 (W0[5:0], PP0[5:0]);
  UB1DCON_6 U25 (W0[6], PP2[6]);
  UB1DCON_7 U26 (W0[7], PP5[7]);
  UB1DCON_8 U27 (W0[8], PP8[8]);
  UB1DCON_14 U28 (W0[14], PP6[14]);
  UB1DCON_15 U29 (W0[15], PP3[15]);
  UBCON_20_16 U30 (W0[20:16], PP0[20:16]);
  UBCON_5_1 U31 (W1[5:1], PP1[5:1]);
  UB1DCON_6 U32 (W1[6], PP3[6]);
  UB1DCON_7 U33 (W1[7], PP6[7]);
  UB1DCON_15 U34 (W1[15], PP4[15]);
  UBCON_19_16 U35 (W1[19:16], PP1[19:16]);
  UBCON_5_2 U36 (W2[5:2], PP2[5:2]);
  UB1DCON_6 U37 (W2[6], PP4[6]);
  UB1DCON_7 U38 (W2[7], PP7[7]);
  UB1DCON_15 U39 (W2[15], PP5[15]);
  UBCON_18_16 U40 (W2[18:16], PP2[18:16]);
  UBCON_5_3 U41 (W3[5:3], PP3[5:3]);
  UB1DCON_6 U42 (W3[6], PP5[6]);
  UBCON_17_16 U43 (W3[17:16], PP3[17:16]);
  UBCON_5_4 U44 (W4[5:4], PP4[5:4]);
  UB1DCON_6 U45 (W4[6], PP6[6]);
  UB1DCON_16 U46 (W4[16], PP4[16]);
  UB1DCON_5 U47 (W5[5], PP5[5]);
  DADTR_20_0_19_1_1001 U48 (S1, S2, W0, W1, W2, W3, W4, W5);
endmodule

module DADTR_20_0_19_1_1001 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5);
  output [20:0] S1;
  output [20:1] S2;
  input [20:0] PP0;
  input [19:1] PP1;
  input [18:2] PP2;
  input [17:3] PP3;
  input [16:4] PP4;
  input [16:5] PP5;
  wire [20:0] W0;
  wire [19:1] W1;
  wire [18:2] W2;
  wire [18:3] W3;
  UBHA_4 U0 (W1[5], W3[4], PP0[4], PP1[4]);
  UBFA_5 U1 (W0[6], W2[5], PP0[5], PP1[5], PP2[5]);
  UBHA_5 U2 (W1[6], W3[5], PP3[5], PP4[5]);
  UBFA_6 U3 (W0[7], W2[6], PP0[6], PP1[6], PP2[6]);
  UBFA_6 U4 (W1[7], W3[6], PP3[6], PP4[6], PP5[6]);
  UBFA_7 U5 (W0[8], W2[7], PP0[7], PP1[7], PP2[7]);
  UBFA_7 U6 (W1[8], W3[7], PP3[7], PP4[7], PP5[7]);
  UBFA_8 U7 (W0[9], W2[8], PP0[8], PP1[8], PP2[8]);
  UBFA_8 U8 (W1[9], W3[8], PP3[8], PP4[8], PP5[8]);
  UBFA_9 U9 (W0[10], W2[9], PP0[9], PP1[9], PP2[9]);
  UBFA_9 U10 (W1[10], W3[9], PP3[9], PP4[9], PP5[9]);
  UBFA_10 U11 (W0[11], W2[10], PP0[10], PP1[10], PP2[10]);
  UBFA_10 U12 (W1[11], W3[10], PP3[10], PP4[10], PP5[10]);
  UBFA_11 U13 (W0[12], W2[11], PP0[11], PP1[11], PP2[11]);
  UBFA_11 U14 (W1[12], W3[11], PP3[11], PP4[11], PP5[11]);
  UBFA_12 U15 (W0[13], W2[12], PP0[12], PP1[12], PP2[12]);
  UBFA_12 U16 (W1[13], W3[12], PP3[12], PP4[12], PP5[12]);
  UBFA_13 U17 (W0[14], W2[13], PP0[13], PP1[13], PP2[13]);
  UBFA_13 U18 (W1[14], W3[13], PP3[13], PP4[13], PP5[13]);
  UBFA_14 U19 (W0[15], W2[14], PP0[14], PP1[14], PP2[14]);
  UBFA_14 U20 (W1[15], W3[14], PP3[14], PP4[14], PP5[14]);
  UBFA_15 U21 (W0[16], W2[15], PP0[15], PP1[15], PP2[15]);
  UBFA_15 U22 (W1[16], W3[15], PP3[15], PP4[15], PP5[15]);
  UBFA_16 U23 (W1[17], W2[16], PP0[16], PP1[16], PP2[16]);
  UBFA_16 U24 (W2[17], W3[16], PP3[16], PP4[16], PP5[16]);
  UBFA_17 U25 (W3[18], W3[17], PP0[17], PP1[17], PP2[17]);
  UBCON_3_0 U26 (W0[3:0], PP0[3:0]);
  UB1DCON_4 U27 (W0[4], PP2[4]);
  UB1DCON_5 U28 (W0[5], PP5[5]);
  UB1DCON_17 U29 (W0[17], PP3[17]);
  UBCON_20_18 U30 (W0[20:18], PP0[20:18]);
  UBCON_3_1 U31 (W1[3:1], PP1[3:1]);
  UB1DCON_4 U32 (W1[4], PP3[4]);
  UBCON_19_18 U33 (W1[19:18], PP1[19:18]);
  UBCON_3_2 U34 (W2[3:2], PP2[3:2]);
  UB1DCON_4 U35 (W2[4], PP4[4]);
  UB1DCON_18 U36 (W2[18], PP2[18]);
  UB1DCON_3 U37 (W3[3], PP3[3]);
  DADTR_20_0_19_1_1002 U38 (S1, S2, W0, W1, W2, W3);
endmodule

module DADTR_20_0_19_1_1002 (S1, S2, PP0, PP1, PP2, PP3);
  output [20:0] S1;
  output [20:1] S2;
  input [20:0] PP0;
  input [19:1] PP1;
  input [18:2] PP2;
  input [18:3] PP3;
  wire [20:0] W0;
  wire [19:1] W1;
  wire [19:2] W2;
  UBHA_3 U0 (W1[4], W2[3], PP0[3], PP1[3]);
  UBFA_4 U1 (W1[5], W2[4], PP0[4], PP1[4], PP2[4]);
  UBFA_5 U2 (W1[6], W2[5], PP0[5], PP1[5], PP2[5]);
  UBFA_6 U3 (W1[7], W2[6], PP0[6], PP1[6], PP2[6]);
  UBFA_7 U4 (W1[8], W2[7], PP0[7], PP1[7], PP2[7]);
  UBFA_8 U5 (W1[9], W2[8], PP0[8], PP1[8], PP2[8]);
  UBFA_9 U6 (W1[10], W2[9], PP0[9], PP1[9], PP2[9]);
  UBFA_10 U7 (W1[11], W2[10], PP0[10], PP1[10], PP2[10]);
  UBFA_11 U8 (W1[12], W2[11], PP0[11], PP1[11], PP2[11]);
  UBFA_12 U9 (W1[13], W2[12], PP0[12], PP1[12], PP2[12]);
  UBFA_13 U10 (W1[14], W2[13], PP0[13], PP1[13], PP2[13]);
  UBFA_14 U11 (W1[15], W2[14], PP0[14], PP1[14], PP2[14]);
  UBFA_15 U12 (W1[16], W2[15], PP0[15], PP1[15], PP2[15]);
  UBFA_16 U13 (W1[17], W2[16], PP0[16], PP1[16], PP2[16]);
  UBFA_17 U14 (W1[18], W2[17], PP0[17], PP1[17], PP2[17]);
  UBFA_18 U15 (W2[19], W2[18], PP0[18], PP1[18], PP2[18]);
  UBCON_2_0 U16 (W0[2:0], PP0[2:0]);
  UB1DCON_3 U17 (W0[3], PP2[3]);
  UBCON_18_4 U18 (W0[18:4], PP3[18:4]);
  UBCON_20_19 U19 (W0[20:19], PP0[20:19]);
  UBCON_2_1 U20 (W1[2:1], PP1[2:1]);
  UB1DCON_3 U21 (W1[3], PP3[3]);
  UB1DCON_19 U22 (W1[19], PP1[19]);
  UB1DCON_2 U23 (W2[2], PP2[2]);
  DADTR_20_0_19_1_1003 U24 (S1, S2, W0, W1, W2);
endmodule

module DADTR_20_0_19_1_1003 (S1, S2, PP0, PP1, PP2);
  output [20:0] S1;
  output [20:1] S2;
  input [20:0] PP0;
  input [19:1] PP1;
  input [19:2] PP2;
  wire [20:0] W0;
  wire [20:1] W1;
  UBHA_2 U0 (W0[3], W1[2], PP0[2], PP1[2]);
  UBFA_3 U1 (W0[4], W1[3], PP0[3], PP1[3], PP2[3]);
  UBFA_4 U2 (W0[5], W1[4], PP0[4], PP1[4], PP2[4]);
  UBFA_5 U3 (W0[6], W1[5], PP0[5], PP1[5], PP2[5]);
  UBFA_6 U4 (W0[7], W1[6], PP0[6], PP1[6], PP2[6]);
  UBFA_7 U5 (W0[8], W1[7], PP0[7], PP1[7], PP2[7]);
  UBFA_8 U6 (W0[9], W1[8], PP0[8], PP1[8], PP2[8]);
  UBFA_9 U7 (W0[10], W1[9], PP0[9], PP1[9], PP2[9]);
  UBFA_10 U8 (W0[11], W1[10], PP0[10], PP1[10], PP2[10]);
  UBFA_11 U9 (W0[12], W1[11], PP0[11], PP1[11], PP2[11]);
  UBFA_12 U10 (W0[13], W1[12], PP0[12], PP1[12], PP2[12]);
  UBFA_13 U11 (W0[14], W1[13], PP0[13], PP1[13], PP2[13]);
  UBFA_14 U12 (W0[15], W1[14], PP0[14], PP1[14], PP2[14]);
  UBFA_15 U13 (W0[16], W1[15], PP0[15], PP1[15], PP2[15]);
  UBFA_16 U14 (W0[17], W1[16], PP0[16], PP1[16], PP2[16]);
  UBFA_17 U15 (W0[18], W1[17], PP0[17], PP1[17], PP2[17]);
  UBFA_18 U16 (W0[19], W1[18], PP0[18], PP1[18], PP2[18]);
  UBFA_19 U17 (W1[20], W1[19], PP0[19], PP1[19], PP2[19]);
  UBCON_1_0 U18 (W0[1:0], PP0[1:0]);
  UB1DCON_2 U19 (W0[2], PP2[2]);
  UB1DCON_20 U20 (W0[20], PP0[20]);
  UB1DCON_1 U21 (W1[1], PP1[1]);
  DADTR_20_0_20_1 U22 (S1, S2, W0, W1);
endmodule

module DADTR_20_0_20_1 (S1, S2, PP0, PP1);
  output [20:0] S1;
  output [20:1] S2;
  input [20:0] PP0;
  input [20:1] PP1;
  UBCON_20_0 U0 (S1, PP0);
  UBCON_20_1 U1 (S2, PP1);
endmodule

module MultUB_STD_DAD_HC000 (P, IN1, IN2);
  output [21:0] P;
  input [11:0] IN1;
  input [9:0] IN2;
  wire [11:0] PP0;
  wire [12:1] PP1;
  wire [13:2] PP2;
  wire [14:3] PP3;
  wire [15:4] PP4;
  wire [16:5] PP5;
  wire [17:6] PP6;
  wire [18:7] PP7;
  wire [19:8] PP8;
  wire [20:9] PP9;
  wire [20:0] S1;
  wire [20:1] S2;
  UBPPG_11_0_9_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, IN1, IN2);
  DADTR_11_0_12_1_1000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9);
  UBHCA_20_0_20_1 U2 (P, S1, S2);
endmodule

module UBCON_12_10 (O, I);
  output [12:10] O;
  input [12:10] I;
  UB1DCON_10 U0 (O[10], I[10]);
  UB1DCON_11 U1 (O[11], I[11]);
  UB1DCON_12 U2 (O[12], I[12]);
endmodule

module UBCON_17_16 (O, I);
  output [17:16] O;
  input [17:16] I;
  UB1DCON_16 U0 (O[16], I[16]);
  UB1DCON_17 U1 (O[17], I[17]);
endmodule

module UBCON_18_16 (O, I);
  output [18:16] O;
  input [18:16] I;
  UB1DCON_16 U0 (O[16], I[16]);
  UB1DCON_17 U1 (O[17], I[17]);
  UB1DCON_18 U2 (O[18], I[18]);
endmodule

module UBCON_18_4 (O, I);
  output [18:4] O;
  input [18:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
  UB1DCON_11 U7 (O[11], I[11]);
  UB1DCON_12 U8 (O[12], I[12]);
  UB1DCON_13 U9 (O[13], I[13]);
  UB1DCON_14 U10 (O[14], I[14]);
  UB1DCON_15 U11 (O[15], I[15]);
  UB1DCON_16 U12 (O[16], I[16]);
  UB1DCON_17 U13 (O[17], I[17]);
  UB1DCON_18 U14 (O[18], I[18]);
endmodule

module UBCON_19_16 (O, I);
  output [19:16] O;
  input [19:16] I;
  UB1DCON_16 U0 (O[16], I[16]);
  UB1DCON_17 U1 (O[17], I[17]);
  UB1DCON_18 U2 (O[18], I[18]);
  UB1DCON_19 U3 (O[19], I[19]);
endmodule

module UBCON_19_18 (O, I);
  output [19:18] O;
  input [19:18] I;
  UB1DCON_18 U0 (O[18], I[18]);
  UB1DCON_19 U1 (O[19], I[19]);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_20_0 (O, I);
  output [20:0] O;
  input [20:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
  UB1DCON_13 U13 (O[13], I[13]);
  UB1DCON_14 U14 (O[14], I[14]);
  UB1DCON_15 U15 (O[15], I[15]);
  UB1DCON_16 U16 (O[16], I[16]);
  UB1DCON_17 U17 (O[17], I[17]);
  UB1DCON_18 U18 (O[18], I[18]);
  UB1DCON_19 U19 (O[19], I[19]);
  UB1DCON_20 U20 (O[20], I[20]);
endmodule

module UBCON_20_1 (O, I);
  output [20:1] O;
  input [20:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
  UB1DCON_6 U5 (O[6], I[6]);
  UB1DCON_7 U6 (O[7], I[7]);
  UB1DCON_8 U7 (O[8], I[8]);
  UB1DCON_9 U8 (O[9], I[9]);
  UB1DCON_10 U9 (O[10], I[10]);
  UB1DCON_11 U10 (O[11], I[11]);
  UB1DCON_12 U11 (O[12], I[12]);
  UB1DCON_13 U12 (O[13], I[13]);
  UB1DCON_14 U13 (O[14], I[14]);
  UB1DCON_15 U14 (O[15], I[15]);
  UB1DCON_16 U15 (O[16], I[16]);
  UB1DCON_17 U16 (O[17], I[17]);
  UB1DCON_18 U17 (O[18], I[18]);
  UB1DCON_19 U18 (O[19], I[19]);
  UB1DCON_20 U19 (O[20], I[20]);
endmodule

module UBCON_20_16 (O, I);
  output [20:16] O;
  input [20:16] I;
  UB1DCON_16 U0 (O[16], I[16]);
  UB1DCON_17 U1 (O[17], I[17]);
  UB1DCON_18 U2 (O[18], I[18]);
  UB1DCON_19 U3 (O[19], I[19]);
  UB1DCON_20 U4 (O[20], I[20]);
endmodule

module UBCON_20_18 (O, I);
  output [20:18] O;
  input [20:18] I;
  UB1DCON_18 U0 (O[18], I[18]);
  UB1DCON_19 U1 (O[19], I[19]);
  UB1DCON_20 U2 (O[20], I[20]);
endmodule

module UBCON_20_19 (O, I);
  output [20:19] O;
  input [20:19] I;
  UB1DCON_19 U0 (O[19], I[19]);
  UB1DCON_20 U1 (O[20], I[20]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBCON_2_1 (O, I);
  output [2:1] O;
  input [2:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
endmodule

module UBCON_3_0 (O, I);
  output [3:0] O;
  input [3:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
endmodule

module UBCON_3_1 (O, I);
  output [3:1] O;
  input [3:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
endmodule

module UBCON_3_2 (O, I);
  output [3:2] O;
  input [3:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
endmodule

module UBCON_5_0 (O, I);
  output [5:0] O;
  input [5:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
endmodule

module UBCON_5_1 (O, I);
  output [5:1] O;
  input [5:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
endmodule

module UBCON_5_2 (O, I);
  output [5:2] O;
  input [5:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
endmodule

module UBCON_5_3 (O, I);
  output [5:3] O;
  input [5:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
endmodule

module UBCON_5_4 (O, I);
  output [5:4] O;
  input [5:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
endmodule

module UBCON_8_0 (O, I);
  output [8:0] O;
  input [8:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
endmodule

module UBCON_8_1 (O, I);
  output [8:1] O;
  input [8:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
  UB1DCON_6 U5 (O[6], I[6]);
  UB1DCON_7 U6 (O[7], I[7]);
  UB1DCON_8 U7 (O[8], I[8]);
endmodule

module UBCON_8_2 (O, I);
  output [8:2] O;
  input [8:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
  UB1DCON_6 U4 (O[6], I[6]);
  UB1DCON_7 U5 (O[7], I[7]);
  UB1DCON_8 U6 (O[8], I[8]);
endmodule

module UBCON_8_3 (O, I);
  output [8:3] O;
  input [8:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
  UB1DCON_6 U3 (O[6], I[6]);
  UB1DCON_7 U4 (O[7], I[7]);
  UB1DCON_8 U5 (O[8], I[8]);
endmodule

module UBCON_8_4 (O, I);
  output [8:4] O;
  input [8:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
endmodule

module UBCON_8_5 (O, I);
  output [8:5] O;
  input [8:5] I;
  UB1DCON_5 U0 (O[5], I[5]);
  UB1DCON_6 U1 (O[6], I[6]);
  UB1DCON_7 U2 (O[7], I[7]);
  UB1DCON_8 U3 (O[8], I[8]);
endmodule

module UBCON_8_6 (O, I);
  output [8:6] O;
  input [8:6] I;
  UB1DCON_6 U0 (O[6], I[6]);
  UB1DCON_7 U1 (O[7], I[7]);
  UB1DCON_8 U2 (O[8], I[8]);
endmodule

module UBCON_8_7 (O, I);
  output [8:7] O;
  input [8:7] I;
  UB1DCON_7 U0 (O[7], I[7]);
  UB1DCON_8 U1 (O[8], I[8]);
endmodule

module UBHCA_20_0_20_1 (S, X, Y);
  output [21:0] S;
  input [20:0] X;
  input [20:1] Y;
  UBPureHCA_20_1 U0 (S[21:1], X[20:1], Y[20:1]);
  UB1DCON_0 U1 (S[0], X[0]);
endmodule

module UBPPG_11_0_9_0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, IN1, IN2);
  output [11:0] PP0;
  output [12:1] PP1;
  output [13:2] PP2;
  output [14:3] PP3;
  output [15:4] PP4;
  output [16:5] PP5;
  output [17:6] PP6;
  output [18:7] PP7;
  output [19:8] PP8;
  output [20:9] PP9;
  input [11:0] IN1;
  input [9:0] IN2;
  UBVPPG_11_0_0 U0 (PP0, IN1, IN2[0]);
  UBVPPG_11_0_1 U1 (PP1, IN1, IN2[1]);
  UBVPPG_11_0_2 U2 (PP2, IN1, IN2[2]);
  UBVPPG_11_0_3 U3 (PP3, IN1, IN2[3]);
  UBVPPG_11_0_4 U4 (PP4, IN1, IN2[4]);
  UBVPPG_11_0_5 U5 (PP5, IN1, IN2[5]);
  UBVPPG_11_0_6 U6 (PP6, IN1, IN2[6]);
  UBVPPG_11_0_7 U7 (PP7, IN1, IN2[7]);
  UBVPPG_11_0_8 U8 (PP8, IN1, IN2[8]);
  UBVPPG_11_0_9 U9 (PP9, IN1, IN2[9]);
endmodule

module UBPureHCA_20_1 (S, X, Y);
  output [21:1] S;
  input [20:1] X;
  input [20:1] Y;
  wire C;
  UBPriHCA_20_1 U0 (S, X, Y, C);
  UBZero_1_1 U1 (C);
endmodule

module UBVPPG_11_0_0 (O, IN1, IN2);
  output [11:0] O;
  input [11:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
  UB1BPPG_6_0 U6 (O[6], IN1[6], IN2);
  UB1BPPG_7_0 U7 (O[7], IN1[7], IN2);
  UB1BPPG_8_0 U8 (O[8], IN1[8], IN2);
  UB1BPPG_9_0 U9 (O[9], IN1[9], IN2);
  UB1BPPG_10_0 U10 (O[10], IN1[10], IN2);
  UB1BPPG_11_0 U11 (O[11], IN1[11], IN2);
endmodule

module UBVPPG_11_0_1 (O, IN1, IN2);
  output [12:1] O;
  input [11:0] IN1;
  input IN2;
  UB1BPPG_0_1 U0 (O[1], IN1[0], IN2);
  UB1BPPG_1_1 U1 (O[2], IN1[1], IN2);
  UB1BPPG_2_1 U2 (O[3], IN1[2], IN2);
  UB1BPPG_3_1 U3 (O[4], IN1[3], IN2);
  UB1BPPG_4_1 U4 (O[5], IN1[4], IN2);
  UB1BPPG_5_1 U5 (O[6], IN1[5], IN2);
  UB1BPPG_6_1 U6 (O[7], IN1[6], IN2);
  UB1BPPG_7_1 U7 (O[8], IN1[7], IN2);
  UB1BPPG_8_1 U8 (O[9], IN1[8], IN2);
  UB1BPPG_9_1 U9 (O[10], IN1[9], IN2);
  UB1BPPG_10_1 U10 (O[11], IN1[10], IN2);
  UB1BPPG_11_1 U11 (O[12], IN1[11], IN2);
endmodule

module UBVPPG_11_0_2 (O, IN1, IN2);
  output [13:2] O;
  input [11:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
  UB1BPPG_6_2 U6 (O[8], IN1[6], IN2);
  UB1BPPG_7_2 U7 (O[9], IN1[7], IN2);
  UB1BPPG_8_2 U8 (O[10], IN1[8], IN2);
  UB1BPPG_9_2 U9 (O[11], IN1[9], IN2);
  UB1BPPG_10_2 U10 (O[12], IN1[10], IN2);
  UB1BPPG_11_2 U11 (O[13], IN1[11], IN2);
endmodule

module UBVPPG_11_0_3 (O, IN1, IN2);
  output [14:3] O;
  input [11:0] IN1;
  input IN2;
  UB1BPPG_0_3 U0 (O[3], IN1[0], IN2);
  UB1BPPG_1_3 U1 (O[4], IN1[1], IN2);
  UB1BPPG_2_3 U2 (O[5], IN1[2], IN2);
  UB1BPPG_3_3 U3 (O[6], IN1[3], IN2);
  UB1BPPG_4_3 U4 (O[7], IN1[4], IN2);
  UB1BPPG_5_3 U5 (O[8], IN1[5], IN2);
  UB1BPPG_6_3 U6 (O[9], IN1[6], IN2);
  UB1BPPG_7_3 U7 (O[10], IN1[7], IN2);
  UB1BPPG_8_3 U8 (O[11], IN1[8], IN2);
  UB1BPPG_9_3 U9 (O[12], IN1[9], IN2);
  UB1BPPG_10_3 U10 (O[13], IN1[10], IN2);
  UB1BPPG_11_3 U11 (O[14], IN1[11], IN2);
endmodule

module UBVPPG_11_0_4 (O, IN1, IN2);
  output [15:4] O;
  input [11:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
  UB1BPPG_6_4 U6 (O[10], IN1[6], IN2);
  UB1BPPG_7_4 U7 (O[11], IN1[7], IN2);
  UB1BPPG_8_4 U8 (O[12], IN1[8], IN2);
  UB1BPPG_9_4 U9 (O[13], IN1[9], IN2);
  UB1BPPG_10_4 U10 (O[14], IN1[10], IN2);
  UB1BPPG_11_4 U11 (O[15], IN1[11], IN2);
endmodule

module UBVPPG_11_0_5 (O, IN1, IN2);
  output [16:5] O;
  input [11:0] IN1;
  input IN2;
  UB1BPPG_0_5 U0 (O[5], IN1[0], IN2);
  UB1BPPG_1_5 U1 (O[6], IN1[1], IN2);
  UB1BPPG_2_5 U2 (O[7], IN1[2], IN2);
  UB1BPPG_3_5 U3 (O[8], IN1[3], IN2);
  UB1BPPG_4_5 U4 (O[9], IN1[4], IN2);
  UB1BPPG_5_5 U5 (O[10], IN1[5], IN2);
  UB1BPPG_6_5 U6 (O[11], IN1[6], IN2);
  UB1BPPG_7_5 U7 (O[12], IN1[7], IN2);
  UB1BPPG_8_5 U8 (O[13], IN1[8], IN2);
  UB1BPPG_9_5 U9 (O[14], IN1[9], IN2);
  UB1BPPG_10_5 U10 (O[15], IN1[10], IN2);
  UB1BPPG_11_5 U11 (O[16], IN1[11], IN2);
endmodule

module UBVPPG_11_0_6 (O, IN1, IN2);
  output [17:6] O;
  input [11:0] IN1;
  input IN2;
  UB1BPPG_0_6 U0 (O[6], IN1[0], IN2);
  UB1BPPG_1_6 U1 (O[7], IN1[1], IN2);
  UB1BPPG_2_6 U2 (O[8], IN1[2], IN2);
  UB1BPPG_3_6 U3 (O[9], IN1[3], IN2);
  UB1BPPG_4_6 U4 (O[10], IN1[4], IN2);
  UB1BPPG_5_6 U5 (O[11], IN1[5], IN2);
  UB1BPPG_6_6 U6 (O[12], IN1[6], IN2);
  UB1BPPG_7_6 U7 (O[13], IN1[7], IN2);
  UB1BPPG_8_6 U8 (O[14], IN1[8], IN2);
  UB1BPPG_9_6 U9 (O[15], IN1[9], IN2);
  UB1BPPG_10_6 U10 (O[16], IN1[10], IN2);
  UB1BPPG_11_6 U11 (O[17], IN1[11], IN2);
endmodule

module UBVPPG_11_0_7 (O, IN1, IN2);
  output [18:7] O;
  input [11:0] IN1;
  input IN2;
  UB1BPPG_0_7 U0 (O[7], IN1[0], IN2);
  UB1BPPG_1_7 U1 (O[8], IN1[1], IN2);
  UB1BPPG_2_7 U2 (O[9], IN1[2], IN2);
  UB1BPPG_3_7 U3 (O[10], IN1[3], IN2);
  UB1BPPG_4_7 U4 (O[11], IN1[4], IN2);
  UB1BPPG_5_7 U5 (O[12], IN1[5], IN2);
  UB1BPPG_6_7 U6 (O[13], IN1[6], IN2);
  UB1BPPG_7_7 U7 (O[14], IN1[7], IN2);
  UB1BPPG_8_7 U8 (O[15], IN1[8], IN2);
  UB1BPPG_9_7 U9 (O[16], IN1[9], IN2);
  UB1BPPG_10_7 U10 (O[17], IN1[10], IN2);
  UB1BPPG_11_7 U11 (O[18], IN1[11], IN2);
endmodule

module UBVPPG_11_0_8 (O, IN1, IN2);
  output [19:8] O;
  input [11:0] IN1;
  input IN2;
  UB1BPPG_0_8 U0 (O[8], IN1[0], IN2);
  UB1BPPG_1_8 U1 (O[9], IN1[1], IN2);
  UB1BPPG_2_8 U2 (O[10], IN1[2], IN2);
  UB1BPPG_3_8 U3 (O[11], IN1[3], IN2);
  UB1BPPG_4_8 U4 (O[12], IN1[4], IN2);
  UB1BPPG_5_8 U5 (O[13], IN1[5], IN2);
  UB1BPPG_6_8 U6 (O[14], IN1[6], IN2);
  UB1BPPG_7_8 U7 (O[15], IN1[7], IN2);
  UB1BPPG_8_8 U8 (O[16], IN1[8], IN2);
  UB1BPPG_9_8 U9 (O[17], IN1[9], IN2);
  UB1BPPG_10_8 U10 (O[18], IN1[10], IN2);
  UB1BPPG_11_8 U11 (O[19], IN1[11], IN2);
endmodule

module UBVPPG_11_0_9 (O, IN1, IN2);
  output [20:9] O;
  input [11:0] IN1;
  input IN2;
  UB1BPPG_0_9 U0 (O[9], IN1[0], IN2);
  UB1BPPG_1_9 U1 (O[10], IN1[1], IN2);
  UB1BPPG_2_9 U2 (O[11], IN1[2], IN2);
  UB1BPPG_3_9 U3 (O[12], IN1[3], IN2);
  UB1BPPG_4_9 U4 (O[13], IN1[4], IN2);
  UB1BPPG_5_9 U5 (O[14], IN1[5], IN2);
  UB1BPPG_6_9 U6 (O[15], IN1[6], IN2);
  UB1BPPG_7_9 U7 (O[16], IN1[7], IN2);
  UB1BPPG_8_9 U8 (O[17], IN1[8], IN2);
  UB1BPPG_9_9 U9 (O[18], IN1[9], IN2);
  UB1BPPG_10_9 U10 (O[19], IN1[10], IN2);
  UB1BPPG_11_9 U11 (O[20], IN1[11], IN2);
endmodule

