/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: Multiplier_6_0_6_000

  Number system: Unsigned binary
  Multiplicand length: 7
  Multiplier length: 7
  Partial product generation: Simple PPG
  Partial product accumulation: Dadda tree
  Final stage addition: Kogge-Stone adder
----------------------------------------------------------------------------*/

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UBHA_6(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_7(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_5(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module GPGenerator(Go, Po, A, B);
  output Go;
  output Po;
  input A;
  input B;
  assign Go = A & B;
  assign Po = A ^ B;
endmodule

module CarryOperator(Go, Po, Gi1, Pi1, Gi2, Pi2);
  output Go;
  output Po;
  input Gi1;
  input Gi2;
  input Pi1;
  input Pi2;
  assign Go = Gi1 | ( Gi2 & Pi1 );
  assign Po = Pi1 & Pi2;
endmodule

module UBPriKSA_12_1(S, X, Y, Cin);
  output [13:1] S;
  input Cin;
  input [12:1] X;
  input [12:1] Y;
  wire [12:1] G0;
  wire [12:1] G1;
  wire [12:1] G2;
  wire [12:1] G3;
  wire [12:1] G4;
  wire [12:1] P0;
  wire [12:1] P1;
  wire [12:1] P2;
  wire [12:1] P3;
  wire [12:1] P4;
  assign P1[1] = P0[1];
  assign G1[1] = G0[1];
  assign P2[1] = P1[1];
  assign G2[1] = G1[1];
  assign P2[2] = P1[2];
  assign G2[2] = G1[2];
  assign P3[1] = P2[1];
  assign G3[1] = G2[1];
  assign P3[2] = P2[2];
  assign G3[2] = G2[2];
  assign P3[3] = P2[3];
  assign G3[3] = G2[3];
  assign P3[4] = P2[4];
  assign G3[4] = G2[4];
  assign P4[1] = P3[1];
  assign G4[1] = G3[1];
  assign P4[2] = P3[2];
  assign G4[2] = G3[2];
  assign P4[3] = P3[3];
  assign G4[3] = G3[3];
  assign P4[4] = P3[4];
  assign G4[4] = G3[4];
  assign P4[5] = P3[5];
  assign G4[5] = G3[5];
  assign P4[6] = P3[6];
  assign G4[6] = G3[6];
  assign P4[7] = P3[7];
  assign G4[7] = G3[7];
  assign P4[8] = P3[8];
  assign G4[8] = G3[8];
  assign S[1] = Cin ^ P0[1];
  assign S[2] = ( G4[1] | ( P4[1] & Cin ) ) ^ P0[2];
  assign S[3] = ( G4[2] | ( P4[2] & Cin ) ) ^ P0[3];
  assign S[4] = ( G4[3] | ( P4[3] & Cin ) ) ^ P0[4];
  assign S[5] = ( G4[4] | ( P4[4] & Cin ) ) ^ P0[5];
  assign S[6] = ( G4[5] | ( P4[5] & Cin ) ) ^ P0[6];
  assign S[7] = ( G4[6] | ( P4[6] & Cin ) ) ^ P0[7];
  assign S[8] = ( G4[7] | ( P4[7] & Cin ) ) ^ P0[8];
  assign S[9] = ( G4[8] | ( P4[8] & Cin ) ) ^ P0[9];
  assign S[10] = ( G4[9] | ( P4[9] & Cin ) ) ^ P0[10];
  assign S[11] = ( G4[10] | ( P4[10] & Cin ) ) ^ P0[11];
  assign S[12] = ( G4[11] | ( P4[11] & Cin ) ) ^ P0[12];
  assign S[13] = G4[12] | ( P4[12] & Cin );
  GPGenerator U0 (G0[1], P0[1], X[1], Y[1]);
  GPGenerator U1 (G0[2], P0[2], X[2], Y[2]);
  GPGenerator U2 (G0[3], P0[3], X[3], Y[3]);
  GPGenerator U3 (G0[4], P0[4], X[4], Y[4]);
  GPGenerator U4 (G0[5], P0[5], X[5], Y[5]);
  GPGenerator U5 (G0[6], P0[6], X[6], Y[6]);
  GPGenerator U6 (G0[7], P0[7], X[7], Y[7]);
  GPGenerator U7 (G0[8], P0[8], X[8], Y[8]);
  GPGenerator U8 (G0[9], P0[9], X[9], Y[9]);
  GPGenerator U9 (G0[10], P0[10], X[10], Y[10]);
  GPGenerator U10 (G0[11], P0[11], X[11], Y[11]);
  GPGenerator U11 (G0[12], P0[12], X[12], Y[12]);
  CarryOperator U12 (G1[2], P1[2], G0[2], P0[2], G0[1], P0[1]);
  CarryOperator U13 (G1[3], P1[3], G0[3], P0[3], G0[2], P0[2]);
  CarryOperator U14 (G1[4], P1[4], G0[4], P0[4], G0[3], P0[3]);
  CarryOperator U15 (G1[5], P1[5], G0[5], P0[5], G0[4], P0[4]);
  CarryOperator U16 (G1[6], P1[6], G0[6], P0[6], G0[5], P0[5]);
  CarryOperator U17 (G1[7], P1[7], G0[7], P0[7], G0[6], P0[6]);
  CarryOperator U18 (G1[8], P1[8], G0[8], P0[8], G0[7], P0[7]);
  CarryOperator U19 (G1[9], P1[9], G0[9], P0[9], G0[8], P0[8]);
  CarryOperator U20 (G1[10], P1[10], G0[10], P0[10], G0[9], P0[9]);
  CarryOperator U21 (G1[11], P1[11], G0[11], P0[11], G0[10], P0[10]);
  CarryOperator U22 (G1[12], P1[12], G0[12], P0[12], G0[11], P0[11]);
  CarryOperator U23 (G2[3], P2[3], G1[3], P1[3], G1[1], P1[1]);
  CarryOperator U24 (G2[4], P2[4], G1[4], P1[4], G1[2], P1[2]);
  CarryOperator U25 (G2[5], P2[5], G1[5], P1[5], G1[3], P1[3]);
  CarryOperator U26 (G2[6], P2[6], G1[6], P1[6], G1[4], P1[4]);
  CarryOperator U27 (G2[7], P2[7], G1[7], P1[7], G1[5], P1[5]);
  CarryOperator U28 (G2[8], P2[8], G1[8], P1[8], G1[6], P1[6]);
  CarryOperator U29 (G2[9], P2[9], G1[9], P1[9], G1[7], P1[7]);
  CarryOperator U30 (G2[10], P2[10], G1[10], P1[10], G1[8], P1[8]);
  CarryOperator U31 (G2[11], P2[11], G1[11], P1[11], G1[9], P1[9]);
  CarryOperator U32 (G2[12], P2[12], G1[12], P1[12], G1[10], P1[10]);
  CarryOperator U33 (G3[5], P3[5], G2[5], P2[5], G2[1], P2[1]);
  CarryOperator U34 (G3[6], P3[6], G2[6], P2[6], G2[2], P2[2]);
  CarryOperator U35 (G3[7], P3[7], G2[7], P2[7], G2[3], P2[3]);
  CarryOperator U36 (G3[8], P3[8], G2[8], P2[8], G2[4], P2[4]);
  CarryOperator U37 (G3[9], P3[9], G2[9], P2[9], G2[5], P2[5]);
  CarryOperator U38 (G3[10], P3[10], G2[10], P2[10], G2[6], P2[6]);
  CarryOperator U39 (G3[11], P3[11], G2[11], P2[11], G2[7], P2[7]);
  CarryOperator U40 (G3[12], P3[12], G2[12], P2[12], G2[8], P2[8]);
  CarryOperator U41 (G4[9], P4[9], G3[9], P3[9], G3[1], P3[1]);
  CarryOperator U42 (G4[10], P4[10], G3[10], P3[10], G3[2], P3[2]);
  CarryOperator U43 (G4[11], P4[11], G3[11], P3[11], G3[3], P3[3]);
  CarryOperator U44 (G4[12], P4[12], G3[12], P3[12], G3[4], P3[4]);
endmodule

module UBZero_1_1(O);
  output [1:1] O;
  assign O[1] = 0;
endmodule

module Multiplier_6_0_6_000(P, IN1, IN2);
  output [13:0] P;
  input [6:0] IN1;
  input [6:0] IN2;
  wire [13:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  assign P[12] = W[12];
  assign P[13] = W[13];
  MultUB_STD_DAD_KS000 U0 (W, IN1, IN2);
endmodule

module DADTR_12_0_11_1_1000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5);
  output [12:0] S1;
  output [12:1] S2;
  input [12:0] PP0;
  input [11:1] PP1;
  input [10:2] PP2;
  input [9:3] PP3;
  input [8:4] PP4;
  input [8:5] PP5;
  wire [12:0] W0;
  wire [11:1] W1;
  wire [10:2] W2;
  wire [10:3] W3;
  UBHA_4 U0 (W1[5], W3[4], PP0[4], PP1[4]);
  UBFA_5 U1 (W0[6], W2[5], PP0[5], PP1[5], PP2[5]);
  UBHA_5 U2 (W1[6], W3[5], PP3[5], PP4[5]);
  UBFA_6 U3 (W0[7], W2[6], PP0[6], PP1[6], PP2[6]);
  UBFA_6 U4 (W1[7], W3[6], PP3[6], PP4[6], PP5[6]);
  UBFA_7 U5 (W0[8], W2[7], PP0[7], PP1[7], PP2[7]);
  UBFA_7 U6 (W1[8], W3[7], PP3[7], PP4[7], PP5[7]);
  UBFA_8 U7 (W1[9], W2[8], PP0[8], PP1[8], PP2[8]);
  UBFA_8 U8 (W2[9], W3[8], PP3[8], PP4[8], PP5[8]);
  UBFA_9 U9 (W3[10], W3[9], PP0[9], PP1[9], PP2[9]);
  UBCON_3_0 U10 (W0[3:0], PP0[3:0]);
  UB1DCON_4 U11 (W0[4], PP2[4]);
  UB1DCON_5 U12 (W0[5], PP5[5]);
  UB1DCON_9 U13 (W0[9], PP3[9]);
  UBCON_12_10 U14 (W0[12:10], PP0[12:10]);
  UBCON_3_1 U15 (W1[3:1], PP1[3:1]);
  UB1DCON_4 U16 (W1[4], PP3[4]);
  UBCON_11_10 U17 (W1[11:10], PP1[11:10]);
  UBCON_3_2 U18 (W2[3:2], PP2[3:2]);
  UB1DCON_4 U19 (W2[4], PP4[4]);
  UB1DCON_10 U20 (W2[10], PP2[10]);
  UB1DCON_3 U21 (W3[3], PP3[3]);
  DADTR_12_0_11_1_1001 U22 (S1, S2, W0, W1, W2, W3);
endmodule

module DADTR_12_0_11_1_1001 (S1, S2, PP0, PP1, PP2, PP3);
  output [12:0] S1;
  output [12:1] S2;
  input [12:0] PP0;
  input [11:1] PP1;
  input [10:2] PP2;
  input [10:3] PP3;
  wire [12:0] W0;
  wire [11:1] W1;
  wire [11:2] W2;
  UBHA_3 U0 (W1[4], W2[3], PP0[3], PP1[3]);
  UBFA_4 U1 (W1[5], W2[4], PP0[4], PP1[4], PP2[4]);
  UBFA_5 U2 (W1[6], W2[5], PP0[5], PP1[5], PP2[5]);
  UBFA_6 U3 (W1[7], W2[6], PP0[6], PP1[6], PP2[6]);
  UBFA_7 U4 (W1[8], W2[7], PP0[7], PP1[7], PP2[7]);
  UBFA_8 U5 (W1[9], W2[8], PP0[8], PP1[8], PP2[8]);
  UBFA_9 U6 (W1[10], W2[9], PP0[9], PP1[9], PP2[9]);
  UBFA_10 U7 (W2[11], W2[10], PP0[10], PP1[10], PP2[10]);
  UBCON_2_0 U8 (W0[2:0], PP0[2:0]);
  UB1DCON_3 U9 (W0[3], PP2[3]);
  UBCON_10_4 U10 (W0[10:4], PP3[10:4]);
  UBCON_12_11 U11 (W0[12:11], PP0[12:11]);
  UBCON_2_1 U12 (W1[2:1], PP1[2:1]);
  UB1DCON_3 U13 (W1[3], PP3[3]);
  UB1DCON_11 U14 (W1[11], PP1[11]);
  UB1DCON_2 U15 (W2[2], PP2[2]);
  DADTR_12_0_11_1_1002 U16 (S1, S2, W0, W1, W2);
endmodule

module DADTR_12_0_11_1_1002 (S1, S2, PP0, PP1, PP2);
  output [12:0] S1;
  output [12:1] S2;
  input [12:0] PP0;
  input [11:1] PP1;
  input [11:2] PP2;
  wire [12:0] W0;
  wire [12:1] W1;
  UBHA_2 U0 (W0[3], W1[2], PP0[2], PP1[2]);
  UBFA_3 U1 (W0[4], W1[3], PP0[3], PP1[3], PP2[3]);
  UBFA_4 U2 (W0[5], W1[4], PP0[4], PP1[4], PP2[4]);
  UBFA_5 U3 (W0[6], W1[5], PP0[5], PP1[5], PP2[5]);
  UBFA_6 U4 (W0[7], W1[6], PP0[6], PP1[6], PP2[6]);
  UBFA_7 U5 (W0[8], W1[7], PP0[7], PP1[7], PP2[7]);
  UBFA_8 U6 (W0[9], W1[8], PP0[8], PP1[8], PP2[8]);
  UBFA_9 U7 (W0[10], W1[9], PP0[9], PP1[9], PP2[9]);
  UBFA_10 U8 (W0[11], W1[10], PP0[10], PP1[10], PP2[10]);
  UBFA_11 U9 (W1[12], W1[11], PP0[11], PP1[11], PP2[11]);
  UBCON_1_0 U10 (W0[1:0], PP0[1:0]);
  UB1DCON_2 U11 (W0[2], PP2[2]);
  UB1DCON_12 U12 (W0[12], PP0[12]);
  UB1DCON_1 U13 (W1[1], PP1[1]);
  DADTR_12_0_12_1 U14 (S1, S2, W0, W1);
endmodule

module DADTR_12_0_12_1 (S1, S2, PP0, PP1);
  output [12:0] S1;
  output [12:1] S2;
  input [12:0] PP0;
  input [12:1] PP1;
  UBCON_12_0 U0 (S1, PP0);
  UBCON_12_1 U1 (S2, PP1);
endmodule

module DADTR_6_0_7_1_8_2000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6);
  output [12:0] S1;
  output [12:1] S2;
  input [6:0] PP0;
  input [7:1] PP1;
  input [8:2] PP2;
  input [9:3] PP3;
  input [10:4] PP4;
  input [11:5] PP5;
  input [12:6] PP6;
  wire [12:0] W0;
  wire [11:1] W1;
  wire [10:2] W2;
  wire [9:3] W3;
  wire [8:4] W4;
  wire [8:5] W5;
  UBHA_6 U0 (W4[7], W5[6], PP0[6], PP1[6]);
  UBHA_7 U1 (W5[8], W5[7], PP1[7], PP2[7]);
  UBCON_5_0 U2 (W0[5:0], PP0[5:0]);
  UB1DCON_6 U3 (W0[6], PP2[6]);
  UB1DCON_7 U4 (W0[7], PP3[7]);
  UB1DCON_8 U5 (W0[8], PP2[8]);
  UB1DCON_9 U6 (W0[9], PP3[9]);
  UB1DCON_10 U7 (W0[10], PP4[10]);
  UB1DCON_11 U8 (W0[11], PP5[11]);
  UB1DCON_12 U9 (W0[12], PP6[12]);
  UBCON_5_1 U10 (W1[5:1], PP1[5:1]);
  UB1DCON_6 U11 (W1[6], PP3[6]);
  UB1DCON_7 U12 (W1[7], PP4[7]);
  UB1DCON_8 U13 (W1[8], PP3[8]);
  UB1DCON_9 U14 (W1[9], PP4[9]);
  UB1DCON_10 U15 (W1[10], PP5[10]);
  UB1DCON_11 U16 (W1[11], PP6[11]);
  UBCON_5_2 U17 (W2[5:2], PP2[5:2]);
  UB1DCON_6 U18 (W2[6], PP4[6]);
  UB1DCON_7 U19 (W2[7], PP5[7]);
  UB1DCON_8 U20 (W2[8], PP4[8]);
  UB1DCON_9 U21 (W2[9], PP5[9]);
  UB1DCON_10 U22 (W2[10], PP6[10]);
  UBCON_5_3 U23 (W3[5:3], PP3[5:3]);
  UB1DCON_6 U24 (W3[6], PP5[6]);
  UB1DCON_7 U25 (W3[7], PP6[7]);
  UB1DCON_8 U26 (W3[8], PP5[8]);
  UB1DCON_9 U27 (W3[9], PP6[9]);
  UBCON_5_4 U28 (W4[5:4], PP4[5:4]);
  UB1DCON_6 U29 (W4[6], PP6[6]);
  UB1DCON_8 U30 (W4[8], PP6[8]);
  UB1DCON_5 U31 (W5[5], PP5[5]);
  DADTR_12_0_11_1_1000 U32 (S1, S2, W0, W1, W2, W3, W4, W5);
endmodule

module MultUB_STD_DAD_KS000 (P, IN1, IN2);
  output [13:0] P;
  input [6:0] IN1;
  input [6:0] IN2;
  wire [6:0] PP0;
  wire [7:1] PP1;
  wire [8:2] PP2;
  wire [9:3] PP3;
  wire [10:4] PP4;
  wire [11:5] PP5;
  wire [12:6] PP6;
  wire [12:0] S1;
  wire [12:1] S2;
  UBPPG_6_0_6_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, IN1, IN2);
  DADTR_6_0_7_1_8_2000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6);
  UBKSA_12_0_12_1 U2 (P, S1, S2);
endmodule

module UBCON_10_4 (O, I);
  output [10:4] O;
  input [10:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
endmodule

module UBCON_11_10 (O, I);
  output [11:10] O;
  input [11:10] I;
  UB1DCON_10 U0 (O[10], I[10]);
  UB1DCON_11 U1 (O[11], I[11]);
endmodule

module UBCON_12_0 (O, I);
  output [12:0] O;
  input [12:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
endmodule

module UBCON_12_1 (O, I);
  output [12:1] O;
  input [12:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
  UB1DCON_6 U5 (O[6], I[6]);
  UB1DCON_7 U6 (O[7], I[7]);
  UB1DCON_8 U7 (O[8], I[8]);
  UB1DCON_9 U8 (O[9], I[9]);
  UB1DCON_10 U9 (O[10], I[10]);
  UB1DCON_11 U10 (O[11], I[11]);
  UB1DCON_12 U11 (O[12], I[12]);
endmodule

module UBCON_12_10 (O, I);
  output [12:10] O;
  input [12:10] I;
  UB1DCON_10 U0 (O[10], I[10]);
  UB1DCON_11 U1 (O[11], I[11]);
  UB1DCON_12 U2 (O[12], I[12]);
endmodule

module UBCON_12_11 (O, I);
  output [12:11] O;
  input [12:11] I;
  UB1DCON_11 U0 (O[11], I[11]);
  UB1DCON_12 U1 (O[12], I[12]);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBCON_2_1 (O, I);
  output [2:1] O;
  input [2:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
endmodule

module UBCON_3_0 (O, I);
  output [3:0] O;
  input [3:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
endmodule

module UBCON_3_1 (O, I);
  output [3:1] O;
  input [3:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
endmodule

module UBCON_3_2 (O, I);
  output [3:2] O;
  input [3:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
endmodule

module UBCON_5_0 (O, I);
  output [5:0] O;
  input [5:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
endmodule

module UBCON_5_1 (O, I);
  output [5:1] O;
  input [5:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
endmodule

module UBCON_5_2 (O, I);
  output [5:2] O;
  input [5:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
endmodule

module UBCON_5_3 (O, I);
  output [5:3] O;
  input [5:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
endmodule

module UBCON_5_4 (O, I);
  output [5:4] O;
  input [5:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
endmodule

module UBKSA_12_0_12_1 (S, X, Y);
  output [13:0] S;
  input [12:0] X;
  input [12:1] Y;
  UBPureKSA_12_1 U0 (S[13:1], X[12:1], Y[12:1]);
  UB1DCON_0 U1 (S[0], X[0]);
endmodule

module UBPPG_6_0_6_0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, IN1, IN2);
  output [6:0] PP0;
  output [7:1] PP1;
  output [8:2] PP2;
  output [9:3] PP3;
  output [10:4] PP4;
  output [11:5] PP5;
  output [12:6] PP6;
  input [6:0] IN1;
  input [6:0] IN2;
  UBVPPG_6_0_0 U0 (PP0, IN1, IN2[0]);
  UBVPPG_6_0_1 U1 (PP1, IN1, IN2[1]);
  UBVPPG_6_0_2 U2 (PP2, IN1, IN2[2]);
  UBVPPG_6_0_3 U3 (PP3, IN1, IN2[3]);
  UBVPPG_6_0_4 U4 (PP4, IN1, IN2[4]);
  UBVPPG_6_0_5 U5 (PP5, IN1, IN2[5]);
  UBVPPG_6_0_6 U6 (PP6, IN1, IN2[6]);
endmodule

module UBPureKSA_12_1 (S, X, Y);
  output [13:1] S;
  input [12:1] X;
  input [12:1] Y;
  wire C;
  UBPriKSA_12_1 U0 (S, X, Y, C);
  UBZero_1_1 U1 (C);
endmodule

module UBVPPG_6_0_0 (O, IN1, IN2);
  output [6:0] O;
  input [6:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
  UB1BPPG_6_0 U6 (O[6], IN1[6], IN2);
endmodule

module UBVPPG_6_0_1 (O, IN1, IN2);
  output [7:1] O;
  input [6:0] IN1;
  input IN2;
  UB1BPPG_0_1 U0 (O[1], IN1[0], IN2);
  UB1BPPG_1_1 U1 (O[2], IN1[1], IN2);
  UB1BPPG_2_1 U2 (O[3], IN1[2], IN2);
  UB1BPPG_3_1 U3 (O[4], IN1[3], IN2);
  UB1BPPG_4_1 U4 (O[5], IN1[4], IN2);
  UB1BPPG_5_1 U5 (O[6], IN1[5], IN2);
  UB1BPPG_6_1 U6 (O[7], IN1[6], IN2);
endmodule

module UBVPPG_6_0_2 (O, IN1, IN2);
  output [8:2] O;
  input [6:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
  UB1BPPG_6_2 U6 (O[8], IN1[6], IN2);
endmodule

module UBVPPG_6_0_3 (O, IN1, IN2);
  output [9:3] O;
  input [6:0] IN1;
  input IN2;
  UB1BPPG_0_3 U0 (O[3], IN1[0], IN2);
  UB1BPPG_1_3 U1 (O[4], IN1[1], IN2);
  UB1BPPG_2_3 U2 (O[5], IN1[2], IN2);
  UB1BPPG_3_3 U3 (O[6], IN1[3], IN2);
  UB1BPPG_4_3 U4 (O[7], IN1[4], IN2);
  UB1BPPG_5_3 U5 (O[8], IN1[5], IN2);
  UB1BPPG_6_3 U6 (O[9], IN1[6], IN2);
endmodule

module UBVPPG_6_0_4 (O, IN1, IN2);
  output [10:4] O;
  input [6:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
  UB1BPPG_6_4 U6 (O[10], IN1[6], IN2);
endmodule

module UBVPPG_6_0_5 (O, IN1, IN2);
  output [11:5] O;
  input [6:0] IN1;
  input IN2;
  UB1BPPG_0_5 U0 (O[5], IN1[0], IN2);
  UB1BPPG_1_5 U1 (O[6], IN1[1], IN2);
  UB1BPPG_2_5 U2 (O[7], IN1[2], IN2);
  UB1BPPG_3_5 U3 (O[8], IN1[3], IN2);
  UB1BPPG_4_5 U4 (O[9], IN1[4], IN2);
  UB1BPPG_5_5 U5 (O[10], IN1[5], IN2);
  UB1BPPG_6_5 U6 (O[11], IN1[6], IN2);
endmodule

module UBVPPG_6_0_6 (O, IN1, IN2);
  output [12:6] O;
  input [6:0] IN1;
  input IN2;
  UB1BPPG_0_6 U0 (O[6], IN1[0], IN2);
  UB1BPPG_1_6 U1 (O[7], IN1[1], IN2);
  UB1BPPG_2_6 U2 (O[8], IN1[2], IN2);
  UB1BPPG_3_6 U3 (O[9], IN1[3], IN2);
  UB1BPPG_4_6 U4 (O[10], IN1[4], IN2);
  UB1BPPG_5_6 U5 (O[11], IN1[5], IN2);
  UB1BPPG_6_6 U6 (O[12], IN1[6], IN2);
endmodule

