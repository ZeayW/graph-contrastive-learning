module CSA_10_0_10_3_11_000 (C, S, X, Y, Z);
  output [11:4] C;
  output [11:0] S;
  input [10:0] X;
  input [10:3] Y;
  input [11:4] Z;
  UBCON_2_0 U0 (S[2:0], X[2:0]);
  UBHA_3 U1 (C[4], S[3], Y[3], X[3]);
  PureCSA_10_4 U2 (C[11:5], S[10:4], Z[10:4], Y[10:4], X[10:4]);
  UB1DCON_11 U3 (S[11], Z[11]);
endmodule

module CSA_11_0_11_4_12_000 (C, S, X, Y, Z);
  output [12:5] C;
  output [12:0] S;
  input [11:0] X;
  input [11:4] Y;
  input [12:5] Z;
  UBCON_3_0 U0 (S[3:0], X[3:0]);
  UBHA_4 U1 (C[5], S[4], Y[4], X[4]);
  PureCSA_11_5 U2 (C[12:6], S[11:5], Z[11:5], Y[11:5], X[11:5]);
  UB1DCON_12 U3 (S[12], Z[12]);
endmodule

module CSA_12_0_12_5_13_000 (C, S, X, Y, Z);
  output [13:6] C;
  output [13:0] S;
  input [12:0] X;
  input [12:5] Y;
  input [13:6] Z;
  UBCON_4_0 U0 (S[4:0], X[4:0]);
  UBHA_5 U1 (C[6], S[5], Y[5], X[5]);
  PureCSA_12_6 U2 (C[13:7], S[12:6], Z[12:6], Y[12:6], X[12:6]);
  UB1DCON_13 U3 (S[13], Z[13]);
endmodule

module CSA_13_0_13_6_14_000 (C, S, X, Y, Z);
  output [14:7] C;
  output [14:0] S;
  input [13:0] X;
  input [13:6] Y;
  input [14:7] Z;
  UBCON_5_0 U0 (S[5:0], X[5:0]);
  UBHA_6 U1 (C[7], S[6], Y[6], X[6]);
  PureCSA_13_7 U2 (C[14:8], S[13:7], Z[13:7], Y[13:7], X[13:7]);
  UB1DCON_14 U3 (S[14], Z[14]);
endmodule

module CSA_7_0_8_1_9_2 (C, S, X, Y, Z);
  output [9:2] C;
  output [9:0] S;
  input [7:0] X;
  input [8:1] Y;
  input [9:2] Z;
  UB1DCON_0 U0 (S[0], X[0]);
  UBHA_1 U1 (C[2], S[1], Y[1], X[1]);
  PureCSA_7_2 U2 (C[8:3], S[7:2], Z[7:2], Y[7:2], X[7:2]);
  UBHA_8 U3 (C[9], S[8], Z[8], Y[8]);
  UB1DCON_9 U4 (S[9], Z[9]);
endmodule

module CSA_9_0_9_2_10_3 (C, S, X, Y, Z);
  output [10:3] C;
  output [10:0] S;
  input [9:0] X;
  input [9:2] Y;
  input [10:3] Z;
  UBCON_1_0 U0 (S[1:0], X[1:0]);
  UBHA_2 U1 (C[3], S[2], Y[2], X[2]);
  PureCSA_9_3 U2 (C[10:4], S[9:3], Z[9:3], Y[9:3], X[9:3]);
  UB1DCON_10 U3 (S[10], Z[10]);
endmodule

module MultUB_STD_ARY_KS000 (P, IN1, IN2);
  output [15:0] P;
  input [7:0] IN1;
  input [7:0] IN2;
  wire [7:0] PP0;
  wire [8:1] PP1;
  wire [9:2] PP2;
  wire [10:3] PP3;
  wire [11:4] PP4;
  wire [12:5] PP5;
  wire [13:6] PP6;
  wire [14:7] PP7;
  wire [14:7] S1;
  wire [14:0] S2;
  UBPPG_7_0_7_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, IN1, IN2);
  UBARYACC_7_0_8_1_000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7);
  UBKSA_14_7_14_0 U2 (P, S1, S2);
endmodule

module PureCSA_10_4 (C, S, X, Y, Z);
  output [11:5] C;
  output [10:4] S;
  input [10:4] X;
  input [10:4] Y;
  input [10:4] Z;
  UBFA_4 U0 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U1 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U2 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U3 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U4 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U5 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U6 (C[11], S[10], X[10], Y[10], Z[10]);
endmodule

module PureCSA_11_5 (C, S, X, Y, Z);
  output [12:6] C;
  output [11:5] S;
  input [11:5] X;
  input [11:5] Y;
  input [11:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U3 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U4 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U5 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U6 (C[12], S[11], X[11], Y[11], Z[11]);
endmodule

module PureCSA_12_6 (C, S, X, Y, Z);
  output [13:7] C;
  output [12:6] S;
  input [12:6] X;
  input [12:6] Y;
  input [12:6] Z;
  UBFA_6 U0 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U1 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U2 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U3 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U4 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U5 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U6 (C[13], S[12], X[12], Y[12], Z[12]);
endmodule

module PureCSA_13_7 (C, S, X, Y, Z);
  output [14:8] C;
  output [13:7] S;
  input [13:7] X;
  input [13:7] Y;
  input [13:7] Z;
  UBFA_7 U0 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U1 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U2 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U3 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U4 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U5 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U6 (C[14], S[13], X[13], Y[13], Z[13]);
endmodule

module PureCSA_7_2 (C, S, X, Y, Z);
  output [8:3] C;
  output [7:2] S;
  input [7:2] X;
  input [7:2] Y;
  input [7:2] Z;
  UBFA_2 U0 (C[3], S[2], X[2], Y[2], Z[2]);
  UBFA_3 U1 (C[4], S[3], X[3], Y[3], Z[3]);
  UBFA_4 U2 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U3 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U4 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U5 (C[8], S[7], X[7], Y[7], Z[7]);
endmodule

module PureCSA_9_3 (C, S, X, Y, Z);
  output [10:4] C;
  output [9:3] S;
  input [9:3] X;
  input [9:3] Y;
  input [9:3] Z;
  UBFA_3 U0 (C[4], S[3], X[3], Y[3], Z[3]);
  UBFA_4 U1 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U2 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U3 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U4 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U5 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U6 (C[10], S[9], X[9], Y[9], Z[9]);
endmodule

module UB1BPPG_0_0 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_0_1 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_0_2 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_0_3 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_0_4 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_0_5 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_0_6 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_0_7 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_1_0 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_1_1 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_1_2 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_1_3 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_1_4 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_1_5 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_1_6 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_1_7 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_2_0 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_2_1 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_2_2 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_2_3 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_2_4 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_2_5 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_2_6 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_2_7 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_3_0 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_3_1 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_3_2 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_3_3 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_3_4 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_3_5 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_3_6 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_3_7 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_4_0 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_4_1 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_4_2 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_4_3 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_4_4 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_4_5 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_4_6 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_4_7 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_5_0 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_5_1 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_5_2 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_5_3 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_5_4 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_5_5 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_5_6 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_5_7 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_6_0 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_6_1 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_6_2 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_6_3 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_6_4 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_6_5 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_6_6 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_6_7 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_7_0 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_7_1 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_7_2 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_7_3 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_7_4 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_7_5 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_7_6 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1BPPG_7_7 (O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
// TODO
endmodule

module UB1DCON_0 (O, I);
  output O;
  input I;
// TODO
endmodule

module UB1DCON_1 (O, I);
  output O;
  input I;
// TODO
endmodule

module UB1DCON_10 (O, I);
  output O;
  input I;
// TODO
endmodule

module UB1DCON_11 (O, I);
  output O;
  input I;
// TODO
endmodule

module UB1DCON_12 (O, I);
  output O;
  input I;
// TODO
endmodule

module UB1DCON_13 (O, I);
  output O;
  input I;
// TODO
endmodule

module UB1DCON_14 (O, I);
  output O;
  input I;
// TODO
endmodule

module UB1DCON_2 (O, I);
  output O;
  input I;
// TODO
endmodule

module UB1DCON_3 (O, I);
  output O;
  input I;
// TODO
endmodule

module UB1DCON_4 (O, I);
  output O;
  input I;
// TODO
endmodule

module UB1DCON_5 (O, I);
  output O;
  input I;
// TODO
endmodule

module UB1DCON_6 (O, I);
  output O;
  input I;
// TODO
endmodule

module UB1DCON_9 (O, I);
  output O;
  input I;
// TODO
endmodule

module UBARYACC_7_0_8_1_000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7);
  output [14:7] S1;
  output [14:0] S2;
  input [7:0] PP0;
  input [8:1] PP1;
  input [9:2] PP2;
  input [10:3] PP3;
  input [11:4] PP4;
  input [12:5] PP5;
  input [13:6] PP6;
  input [14:7] PP7;
  wire [9:2] IC0;
  wire [10:3] IC1;
  wire [11:4] IC2;
  wire [12:5] IC3;
  wire [13:6] IC4;
  wire [9:0] IS0;
  wire [10:0] IS1;
  wire [11:0] IS2;
  wire [12:0] IS3;
  wire [13:0] IS4;
  CSA_7_0_8_1_9_2 U0 (IC0, IS0, PP0, PP1, PP2);
  CSA_9_0_9_2_10_3 U1 (IC1, IS1, IS0, IC0, PP3);
  CSA_10_0_10_3_11_000 U2 (IC2, IS2, IS1, IC1, PP4);
  CSA_11_0_11_4_12_000 U3 (IC3, IS3, IS2, IC2, PP5);
  CSA_12_0_12_5_13_000 U4 (IC4, IS4, IS3, IC3, PP6);
  CSA_13_0_13_6_14_000 U5 (S1, S2, IS4, IC4, PP7);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBCON_3_0 (O, I);
  output [3:0] O;
  input [3:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
endmodule

module UBCON_4_0 (O, I);
  output [4:0] O;
  input [4:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
endmodule

module UBCON_5_0 (O, I);
  output [5:0] O;
  input [5:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
endmodule

module UBCON_6_0 (O, I);
  output [6:0] O;
  input [6:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
endmodule

module UBFA_10 (C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
// TODO
endmodule

module UBFA_11 (C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
// TODO
endmodule

module UBFA_12 (C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
// TODO
endmodule

module UBFA_13 (C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
// TODO
endmodule

module UBFA_2 (C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
// TODO
endmodule

module UBFA_3 (C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
// TODO
endmodule

module UBFA_4 (C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
// TODO
endmodule

module UBFA_5 (C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
// TODO
endmodule

module UBFA_6 (C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
// TODO
endmodule

module UBFA_7 (C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
// TODO
endmodule

module UBFA_8 (C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
// TODO
endmodule

module UBFA_9 (C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
// TODO
endmodule

module UBHA_1 (C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
// TODO
endmodule

module UBHA_2 (C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
// TODO
endmodule

module UBHA_3 (C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
// TODO
endmodule

module UBHA_4 (C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
// TODO
endmodule

module UBHA_5 (C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
// TODO
endmodule

module UBHA_6 (C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
// TODO
endmodule

module UBHA_8 (C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
// TODO
endmodule

module UBKSA_14_7_14_0 (S, X, Y);
  output [15:0] S;
  input [14:7] X;
  input [14:0] Y;
  UBPureKSA_14_7 U0 (S[15:7], X[14:7], Y[14:7]);
  UBCON_6_0 U1 (S[6:0], Y[6:0]);
endmodule

module UBPPG_7_0_7_0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, IN1, IN2);
  output [7:0] PP0;
  output [8:1] PP1;
  output [9:2] PP2;
  output [10:3] PP3;
  output [11:4] PP4;
  output [12:5] PP5;
  output [13:6] PP6;
  output [14:7] PP7;
  input [7:0] IN1;
  input [7:0] IN2;
  UBVPPG_7_0_0 U0 (PP0, IN1, IN2[0]);
  UBVPPG_7_0_1 U1 (PP1, IN1, IN2[1]);
  UBVPPG_7_0_2 U2 (PP2, IN1, IN2[2]);
  UBVPPG_7_0_3 U3 (PP3, IN1, IN2[3]);
  UBVPPG_7_0_4 U4 (PP4, IN1, IN2[4]);
  UBVPPG_7_0_5 U5 (PP5, IN1, IN2[5]);
  UBVPPG_7_0_6 U6 (PP6, IN1, IN2[6]);
  UBVPPG_7_0_7 U7 (PP7, IN1, IN2[7]);
endmodule

module UBPriKSA_14_7 (S, X, Y, Cin);
  output [15:7] S;
  input Cin;
  input [14:7] X;
  input [14:7] Y;
// TODO
endmodule

module UBPureKSA_14_7 (S, X, Y);
  output [15:7] S;
  input [14:7] X;
  input [14:7] Y;
  wire C;
  UBPriKSA_14_7 U0 (S, X, Y, C);
  UBZero_7_7 U1 (C);
endmodule

module UBVPPG_7_0_0 (O, IN1, IN2);
  output [7:0] O;
  input [7:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
  UB1BPPG_6_0 U6 (O[6], IN1[6], IN2);
  UB1BPPG_7_0 U7 (O[7], IN1[7], IN2);
endmodule

module UBVPPG_7_0_1 (O, IN1, IN2);
  output [8:1] O;
  input [7:0] IN1;
  input IN2;
  UB1BPPG_0_1 U0 (O[1], IN1[0], IN2);
  UB1BPPG_1_1 U1 (O[2], IN1[1], IN2);
  UB1BPPG_2_1 U2 (O[3], IN1[2], IN2);
  UB1BPPG_3_1 U3 (O[4], IN1[3], IN2);
  UB1BPPG_4_1 U4 (O[5], IN1[4], IN2);
  UB1BPPG_5_1 U5 (O[6], IN1[5], IN2);
  UB1BPPG_6_1 U6 (O[7], IN1[6], IN2);
  UB1BPPG_7_1 U7 (O[8], IN1[7], IN2);
endmodule

module UBVPPG_7_0_2 (O, IN1, IN2);
  output [9:2] O;
  input [7:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
  UB1BPPG_6_2 U6 (O[8], IN1[6], IN2);
  UB1BPPG_7_2 U7 (O[9], IN1[7], IN2);
endmodule

module UBVPPG_7_0_3 (O, IN1, IN2);
  output [10:3] O;
  input [7:0] IN1;
  input IN2;
  UB1BPPG_0_3 U0 (O[3], IN1[0], IN2);
  UB1BPPG_1_3 U1 (O[4], IN1[1], IN2);
  UB1BPPG_2_3 U2 (O[5], IN1[2], IN2);
  UB1BPPG_3_3 U3 (O[6], IN1[3], IN2);
  UB1BPPG_4_3 U4 (O[7], IN1[4], IN2);
  UB1BPPG_5_3 U5 (O[8], IN1[5], IN2);
  UB1BPPG_6_3 U6 (O[9], IN1[6], IN2);
  UB1BPPG_7_3 U7 (O[10], IN1[7], IN2);
endmodule

module UBVPPG_7_0_4 (O, IN1, IN2);
  output [11:4] O;
  input [7:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
  UB1BPPG_6_4 U6 (O[10], IN1[6], IN2);
  UB1BPPG_7_4 U7 (O[11], IN1[7], IN2);
endmodule

module UBVPPG_7_0_5 (O, IN1, IN2);
  output [12:5] O;
  input [7:0] IN1;
  input IN2;
  UB1BPPG_0_5 U0 (O[5], IN1[0], IN2);
  UB1BPPG_1_5 U1 (O[6], IN1[1], IN2);
  UB1BPPG_2_5 U2 (O[7], IN1[2], IN2);
  UB1BPPG_3_5 U3 (O[8], IN1[3], IN2);
  UB1BPPG_4_5 U4 (O[9], IN1[4], IN2);
  UB1BPPG_5_5 U5 (O[10], IN1[5], IN2);
  UB1BPPG_6_5 U6 (O[11], IN1[6], IN2);
  UB1BPPG_7_5 U7 (O[12], IN1[7], IN2);
endmodule

module UBVPPG_7_0_6 (O, IN1, IN2);
  output [13:6] O;
  input [7:0] IN1;
  input IN2;
  UB1BPPG_0_6 U0 (O[6], IN1[0], IN2);
  UB1BPPG_1_6 U1 (O[7], IN1[1], IN2);
  UB1BPPG_2_6 U2 (O[8], IN1[2], IN2);
  UB1BPPG_3_6 U3 (O[9], IN1[3], IN2);
  UB1BPPG_4_6 U4 (O[10], IN1[4], IN2);
  UB1BPPG_5_6 U5 (O[11], IN1[5], IN2);
  UB1BPPG_6_6 U6 (O[12], IN1[6], IN2);
  UB1BPPG_7_6 U7 (O[13], IN1[7], IN2);
endmodule

module UBVPPG_7_0_7 (O, IN1, IN2);
  output [14:7] O;
  input [7:0] IN1;
  input IN2;
  UB1BPPG_0_7 U0 (O[7], IN1[0], IN2);
  UB1BPPG_1_7 U1 (O[8], IN1[1], IN2);
  UB1BPPG_2_7 U2 (O[9], IN1[2], IN2);
  UB1BPPG_3_7 U3 (O[10], IN1[3], IN2);
  UB1BPPG_4_7 U4 (O[11], IN1[4], IN2);
  UB1BPPG_5_7 U5 (O[12], IN1[5], IN2);
  UB1BPPG_6_7 U6 (O[13], IN1[6], IN2);
  UB1BPPG_7_7 U7 (O[14], IN1[7], IN2);
endmodule

module UBZero_7_7 (O);
  output O;
// TODO
endmodule

