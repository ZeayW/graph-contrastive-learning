/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: UBCLA_30_0_30_0

  Operand-1 length: 31
  Operand-2 length: 31
  Two-operand addition algorithm: Carry look-ahead adder
----------------------------------------------------------------------------*/

module GPGenerator(Go, Po, A, B);
  output Go;
  output Po;
  input A;
  input B;
  assign Go = A & B;
  assign Po = A ^ B;
endmodule

module CLAUnit_31(C, G, P, Cin);
  output [31:1] C;
  input Cin;
  input [30:0] G;
  input [30:0] P;
  assign C[1] = G[0] | ( P[0] & Cin );
  assign C[2] = G[1] | ( P[1] & G[0] ) | ( P[1] & P[0] & Cin );
  assign C[3] = G[2] | ( P[2] & G[1] ) | ( P[2] & P[1] & G[0] ) | ( P[2] & P[1] & P[0] & Cin );
  assign C[4] = G[3] | ( P[3] & G[2] ) | ( P[3] & P[2] & G[1] ) | ( P[3] & P[2] & P[1] & G[0] ) | ( P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[5] = G[4] | ( P[4] & G[3] ) | ( P[4] & P[3] & G[2] ) | ( P[4] & P[3] & P[2] & G[1] ) | ( P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[6] = G[5] | ( P[5] & G[4] ) | ( P[5] & P[4] & G[3] ) | ( P[5] & P[4] & P[3] & G[2] ) | ( P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[5] & P[4] & P[3]
 & P[2] & P[1] & P[0] & Cin );
  assign C[7] = G[6] | ( P[6] & G[5] ) | ( P[6] & P[5] & G[4] ) | ( P[6] & P[5] & P[4] & G[3] ) | ( P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[6] & P[5] & P[4]
 & P[3] & P[2] & P[1] & G[0] ) | ( P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[8] = G[7] | ( P[7] & G[6] ) | ( P[7] & P[6] & G[5] ) | ( P[7] & P[6] & P[5] & G[4] ) | ( P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[7] & P[6] & P[5]
 & P[4] & P[3] & P[2] & G[1] ) | ( P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[9] = G[8] | ( P[8] & G[7] ) | ( P[8] & P[7] & G[6] ) | ( P[8] & P[7] & P[6] & G[5] ) | ( P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & G[2] ) | ( P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[8] & P[7] & P[6] & P[5] & P[4] & P[3]
 & P[2] & P[1] & P[0] & Cin );
  assign C[10] = G[9] | ( P[9] & G[8] ) | ( P[9] & P[8] & G[7] ) | ( P[9] & P[8] & P[7] & G[6] ) | ( P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & G[3] ) | ( P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & P[1] & G[0] ) | ( P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[11] = G[10] | ( P[10] & G[9] ) | ( P[10] & P[9] & G[8] ) | ( P[10] & P[9] & P[8] & G[7] ) | ( P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] &
 Cin );
  assign C[12] = G[11] | ( P[11] & G[10] ) | ( P[11] & P[10] & G[9] ) | ( P[11] & P[10] & P[9] & G[8] ) | ( P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[11]
 & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[11] & P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3]
 & P[2] & P[1] & G[0] ) | ( P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[13] = G[12] | ( P[12] & G[11] ) | ( P[12] & P[11] & G[10] ) | ( P[12] & P[11] & P[10] & G[9] ) | ( P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & G[1] ) | ( P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2]
 & P[1] & P[0] & Cin );
  assign C[14] = G[13] | ( P[13] & G[12] ) | ( P[13] & P[12] & G[11] ) | ( P[13] & P[12] & P[11] & G[10] ) | ( P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) |
 ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[13] &
 P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] &
 P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[15] = G[14] | ( P[14] & G[13] ) | ( P[14] & P[13] & G[12] ) | ( P[14] & P[13] & P[12] & G[11] ) | ( P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & G[9] )
 | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] &
 P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[16] = G[15] | ( P[15] & G[14] ) | ( P[15] & P[14] & G[13] ) | ( P[15] & P[14] & P[13] & G[12] ) | ( P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & G[10] )
 | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | (
 P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[15] & P[14] & P[13] &
 P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] &
 P[1] & P[0] & Cin );
  assign C[17] = G[16] | ( P[16] & G[15] ) | ( P[16] & P[15] & G[14] ) | ( P[16] & P[15] & P[14] & G[13] ) | ( P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & G[11] )
 | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] )
 | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[16] & P[15]
 & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & P[1] & G[0] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[18] = G[17] | ( P[17] & G[16] ) | ( P[17] & P[16] & G[15] ) | ( P[17] & P[16] & P[15] & G[14] ) | ( P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & G[12] )
 | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9]
 ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[17] & P[16] &
 P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[19] = G[18] | ( P[18] & G[17] ) | ( P[18] & P[17] & G[16] ) | ( P[18] & P[17] & P[16] & G[15] ) | ( P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & G[13] )
 | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10]
 ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4]
 ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | (
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] &
 P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[20] = G[19] | ( P[19] & G[18] ) | ( P[19] & P[18] & G[17] ) | ( P[19] & P[18] & P[17] & G[16] ) | ( P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & G[14] )
 | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11]
 ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5]
 ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) |
 ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] &
 P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[21] = G[20] | ( P[20] & G[19] ) | ( P[20] & P[19] & G[18] ) | ( P[20] & P[19] & P[18] & G[17] ) | ( P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & G[15] )
 | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12]
 ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6]
 ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] )
 | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8]
 & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2]
 & P[1] & P[0] & Cin );
  assign C[22] = G[21] | ( P[21] & G[20] ) | ( P[21] & P[20] & G[19] ) | ( P[21] & P[20] & P[19] & G[18] ) | ( P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & G[16] )
 | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13]
 ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[21] & P[20] & P[19]
 & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] &
 P[8] & G[7] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & G[4] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] &
 P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2]
 & P[1] & P[0] & Cin );
  assign C[23] = G[22] | ( P[22] & G[21] ) | ( P[22] & P[21] & G[20] ) | ( P[22] & P[21] & P[20] & G[19] ) | ( P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & G[17] )
 | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14]
 ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & G[8] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & G[5] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8]
 & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] &
 P[3] & P[2] & P[1] & G[0] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0]
 & Cin );
  assign C[24] = G[23] | ( P[23] & G[22] ) | ( P[23] & P[22] & G[21] ) | ( P[23] & P[22] & P[21] & G[20] ) | ( P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & G[18] )
 | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15]
 ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & G[9] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] &
 P[8] & P[7] & G[6] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] &
 P[4] & P[3] & P[2] & G[1] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1]
 & G[0] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[25] = G[24] | ( P[24] & G[23] ) | ( P[24] & P[23] & G[22] ) | ( P[24] & P[23] & P[22] & G[21] ) | ( P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & G[19] )
 | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16]
 ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & G[10] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] &
 P[10] & P[9] & P[8] & G[7] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8]
 & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5]
 & P[4] & P[3] & P[2] & G[1] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3]
 & P[2] & P[1] & G[0] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2]
 & P[1] & P[0] & Cin );
  assign C[26] = G[25] | ( P[25] & G[24] ) | ( P[25] & P[24] & G[23] ) | ( P[25] & P[24] & P[23] & G[22] ) | ( P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & G[20] )
 | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17]
 ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & G[11] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & G[8] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5]
 & P[4] & P[3] & P[2] & G[1] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & P[1] & G[0] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[27] = G[26] | ( P[26] & G[25] ) | ( P[26] & P[25] & G[24] ) | ( P[26] & P[25] & P[24] & G[23] ) | ( P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & G[21] )
 | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18]
 ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[26] & P[25] &
 P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & G[12] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & G[9] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] &
 P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[28] = G[27] | ( P[27] & G[26] ) | ( P[27] & P[26] & G[25] ) | ( P[27] & P[26] & P[25] & G[24] ) | ( P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & G[22] )
 | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19]
 ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[27] & P[26] &
 P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & G[13] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & G[10] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] &
 P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[29] = G[28] | ( P[28] & G[27] ) | ( P[28] & P[27] & G[26] ) | ( P[28] & P[27] & P[26] & G[25] ) | ( P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & G[23] )
 | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20]
 ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & G[14] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & P[13] & P[12] & G[11] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19]
 & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[30] = G[29] | ( P[29] & G[28] ) | ( P[29] & P[28] & G[27] ) | ( P[29] & P[28] & P[27] & G[26] ) | ( P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & G[24] )
 | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21]
 ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[29] & P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & G[15] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & G[12] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19]
 & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[31] = G[30] | ( P[30] & G[29] ) | ( P[30] & P[29] & G[28] ) | ( P[30] & P[29] & P[28] & G[27] ) | ( P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & G[25] )
 | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22]
 ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & G[16] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] &
 P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & G[13] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[30] &
 P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & P[1] & P[0] & Cin );
endmodule

module UBPriCLA_30_0(S, X, Y, Cin);
  output [31:0] S;
  input Cin;
  input [30:0] X;
  input [30:0] Y;
  wire [31:1] C;
  wire [30:0] G;
  wire [30:0] P;
  assign S[0] = Cin ^ P[0];
  assign S[1] = C[1] ^ P[1];
  assign S[2] = C[2] ^ P[2];
  assign S[3] = C[3] ^ P[3];
  assign S[4] = C[4] ^ P[4];
  assign S[5] = C[5] ^ P[5];
  assign S[6] = C[6] ^ P[6];
  assign S[7] = C[7] ^ P[7];
  assign S[8] = C[8] ^ P[8];
  assign S[9] = C[9] ^ P[9];
  assign S[10] = C[10] ^ P[10];
  assign S[11] = C[11] ^ P[11];
  assign S[12] = C[12] ^ P[12];
  assign S[13] = C[13] ^ P[13];
  assign S[14] = C[14] ^ P[14];
  assign S[15] = C[15] ^ P[15];
  assign S[16] = C[16] ^ P[16];
  assign S[17] = C[17] ^ P[17];
  assign S[18] = C[18] ^ P[18];
  assign S[19] = C[19] ^ P[19];
  assign S[20] = C[20] ^ P[20];
  assign S[21] = C[21] ^ P[21];
  assign S[22] = C[22] ^ P[22];
  assign S[23] = C[23] ^ P[23];
  assign S[24] = C[24] ^ P[24];
  assign S[25] = C[25] ^ P[25];
  assign S[26] = C[26] ^ P[26];
  assign S[27] = C[27] ^ P[27];
  assign S[28] = C[28] ^ P[28];
  assign S[29] = C[29] ^ P[29];
  assign S[30] = C[30] ^ P[30];
  assign S[31] = C[31];
  GPGenerator U0 (G[0], P[0], X[0], Y[0]);
  GPGenerator U1 (G[1], P[1], X[1], Y[1]);
  GPGenerator U2 (G[2], P[2], X[2], Y[2]);
  GPGenerator U3 (G[3], P[3], X[3], Y[3]);
  GPGenerator U4 (G[4], P[4], X[4], Y[4]);
  GPGenerator U5 (G[5], P[5], X[5], Y[5]);
  GPGenerator U6 (G[6], P[6], X[6], Y[6]);
  GPGenerator U7 (G[7], P[7], X[7], Y[7]);
  GPGenerator U8 (G[8], P[8], X[8], Y[8]);
  GPGenerator U9 (G[9], P[9], X[9], Y[9]);
  GPGenerator U10 (G[10], P[10], X[10], Y[10]);
  GPGenerator U11 (G[11], P[11], X[11], Y[11]);
  GPGenerator U12 (G[12], P[12], X[12], Y[12]);
  GPGenerator U13 (G[13], P[13], X[13], Y[13]);
  GPGenerator U14 (G[14], P[14], X[14], Y[14]);
  GPGenerator U15 (G[15], P[15], X[15], Y[15]);
  GPGenerator U16 (G[16], P[16], X[16], Y[16]);
  GPGenerator U17 (G[17], P[17], X[17], Y[17]);
  GPGenerator U18 (G[18], P[18], X[18], Y[18]);
  GPGenerator U19 (G[19], P[19], X[19], Y[19]);
  GPGenerator U20 (G[20], P[20], X[20], Y[20]);
  GPGenerator U21 (G[21], P[21], X[21], Y[21]);
  GPGenerator U22 (G[22], P[22], X[22], Y[22]);
  GPGenerator U23 (G[23], P[23], X[23], Y[23]);
  GPGenerator U24 (G[24], P[24], X[24], Y[24]);
  GPGenerator U25 (G[25], P[25], X[25], Y[25]);
  GPGenerator U26 (G[26], P[26], X[26], Y[26]);
  GPGenerator U27 (G[27], P[27], X[27], Y[27]);
  GPGenerator U28 (G[28], P[28], X[28], Y[28]);
  GPGenerator U29 (G[29], P[29], X[29], Y[29]);
  GPGenerator U30 (G[30], P[30], X[30], Y[30]);
  CLAUnit_31 U31 (C, G, P, Cin);
endmodule

module UBZero_0_0(O);
  output [0:0] O;
  assign O[0] = 0;
endmodule

module UBCLA_30_0_30_0 (S, X, Y);
  output [31:0] S;
  input [30:0] X;
  input [30:0] Y;
  UBPureCLA_30_0 U0 (S[31:0], X[30:0], Y[30:0]);
endmodule

module UBPureCLA_30_0 (S, X, Y);
  output [31:0] S;
  input [30:0] X;
  input [30:0] Y;
  wire C;
  UBPriCLA_30_0 U0 (S, X, Y, C);
  UBZero_0_0 U1 (C);
endmodule

