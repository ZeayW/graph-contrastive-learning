/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: Multiplier_13_0_1000

  Number system: Unsigned binary
  Multiplicand length: 14
  Multiplier length: 14
  Partial product generation: Simple PPG
  Partial product accumulation: (7,3) counter tree
  Final stage addition: Kogge-Stone adder
----------------------------------------------------------------------------*/

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UBHA_7(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB4_3C8(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C9(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C10(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C11(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBHA_11(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB7_3C12(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C12(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C13(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C13(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C14(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C14(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C15(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C15(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C16(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_16(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB7_3C17(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBHA_17(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB6_3C18(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C19(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_20(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_21(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_21(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_23(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_24(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_25(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB4_3C4(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB5_3C5(S1, S2, S3, X1, X2, X3, X4, X5);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = X4 & X5;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C6(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C7(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C8(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C9(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C18(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C19(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C20(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB7_3C21(S1, S2, S3, X1, X2, X3, X4, X5, X6, X7);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  input X7;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 ^ X7 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & ( X6 | X7 ) ) ) & ( ~ ( ( X4 & X5 ) | ( X6 & X7 ) ) ) );
  assign W5 = ~ ( X4 & X5 & X6 & X7 );
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB6_3C22(S1, S2, S3, X1, X2, X3, X4, X5, X6);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  input X5;
  input X6;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4 ^ X5 ^ ( X6 );
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = ~ ( ( ~ ( ( X4 | X5 ) & X6 ) ) & ( ~ ( X4 & X5 ) ) );
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UB4_3C23(S1, S2, S3, X1, X2, X3, X4);
  output S1;
  output S2;
  output S3;
  input X1;
  input X2;
  input X3;
  input X4;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  assign W1 = X1 ^ X2 ^ X3;
  assign W2 = X4;
  assign W3 = ~ ( ( ~ ( X1 & X2 ) ) & ( ~ ( X1 & X3 ) ) & ( ~ ( X2 & X3 ) ) );
  assign W4 = 0;
  assign W5 = 1;
  assign W6 = ~ ( ( ~ ( W4 & W5 ) ) ^ W3 );
  assign S3 = W1 ^ W2;
  assign S2 = ~ ( W6 ^ ( ~ ( W1 & W2 ) ) );
  assign S1 = ~ ( W5 & ( ~ ( W3 & W4 ) ) & ( ~ ( W1 & W2 & W6 ) ) );
endmodule

module UBFA_24(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_25(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_12(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_13(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_14(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_15(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_17(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_18(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_19(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_21(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_22(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_23(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_25(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_26(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_27(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_27_27(O);
  output [27:27] O;
  assign O[27] = 0;
endmodule

module GPGenerator(Go, Po, A, B);
  output Go;
  output Po;
  input A;
  input B;
  assign Go = A & B;
  assign Po = A ^ B;
endmodule

module CarryOperator(Go, Po, Gi1, Pi1, Gi2, Pi2);
  output Go;
  output Po;
  input Gi1;
  input Gi2;
  input Pi1;
  input Pi2;
  assign Go = Gi1 | ( Gi2 & Pi1 );
  assign Po = Pi1 & Pi2;
endmodule

module UBPriKSA_27_1(S, X, Y, Cin);
  output [28:1] S;
  input Cin;
  input [27:1] X;
  input [27:1] Y;
  wire [27:1] G0;
  wire [27:1] G1;
  wire [27:1] G2;
  wire [27:1] G3;
  wire [27:1] G4;
  wire [27:1] G5;
  wire [27:1] P0;
  wire [27:1] P1;
  wire [27:1] P2;
  wire [27:1] P3;
  wire [27:1] P4;
  wire [27:1] P5;
  assign P1[1] = P0[1];
  assign G1[1] = G0[1];
  assign P2[1] = P1[1];
  assign G2[1] = G1[1];
  assign P2[2] = P1[2];
  assign G2[2] = G1[2];
  assign P3[1] = P2[1];
  assign G3[1] = G2[1];
  assign P3[2] = P2[2];
  assign G3[2] = G2[2];
  assign P3[3] = P2[3];
  assign G3[3] = G2[3];
  assign P3[4] = P2[4];
  assign G3[4] = G2[4];
  assign P4[1] = P3[1];
  assign G4[1] = G3[1];
  assign P4[2] = P3[2];
  assign G4[2] = G3[2];
  assign P4[3] = P3[3];
  assign G4[3] = G3[3];
  assign P4[4] = P3[4];
  assign G4[4] = G3[4];
  assign P4[5] = P3[5];
  assign G4[5] = G3[5];
  assign P4[6] = P3[6];
  assign G4[6] = G3[6];
  assign P4[7] = P3[7];
  assign G4[7] = G3[7];
  assign P4[8] = P3[8];
  assign G4[8] = G3[8];
  assign P5[1] = P4[1];
  assign G5[1] = G4[1];
  assign P5[2] = P4[2];
  assign G5[2] = G4[2];
  assign P5[3] = P4[3];
  assign G5[3] = G4[3];
  assign P5[4] = P4[4];
  assign G5[4] = G4[4];
  assign P5[5] = P4[5];
  assign G5[5] = G4[5];
  assign P5[6] = P4[6];
  assign G5[6] = G4[6];
  assign P5[7] = P4[7];
  assign G5[7] = G4[7];
  assign P5[8] = P4[8];
  assign G5[8] = G4[8];
  assign P5[9] = P4[9];
  assign G5[9] = G4[9];
  assign P5[10] = P4[10];
  assign G5[10] = G4[10];
  assign P5[11] = P4[11];
  assign G5[11] = G4[11];
  assign P5[12] = P4[12];
  assign G5[12] = G4[12];
  assign P5[13] = P4[13];
  assign G5[13] = G4[13];
  assign P5[14] = P4[14];
  assign G5[14] = G4[14];
  assign P5[15] = P4[15];
  assign G5[15] = G4[15];
  assign P5[16] = P4[16];
  assign G5[16] = G4[16];
  assign S[1] = Cin ^ P0[1];
  assign S[2] = ( G5[1] | ( P5[1] & Cin ) ) ^ P0[2];
  assign S[3] = ( G5[2] | ( P5[2] & Cin ) ) ^ P0[3];
  assign S[4] = ( G5[3] | ( P5[3] & Cin ) ) ^ P0[4];
  assign S[5] = ( G5[4] | ( P5[4] & Cin ) ) ^ P0[5];
  assign S[6] = ( G5[5] | ( P5[5] & Cin ) ) ^ P0[6];
  assign S[7] = ( G5[6] | ( P5[6] & Cin ) ) ^ P0[7];
  assign S[8] = ( G5[7] | ( P5[7] & Cin ) ) ^ P0[8];
  assign S[9] = ( G5[8] | ( P5[8] & Cin ) ) ^ P0[9];
  assign S[10] = ( G5[9] | ( P5[9] & Cin ) ) ^ P0[10];
  assign S[11] = ( G5[10] | ( P5[10] & Cin ) ) ^ P0[11];
  assign S[12] = ( G5[11] | ( P5[11] & Cin ) ) ^ P0[12];
  assign S[13] = ( G5[12] | ( P5[12] & Cin ) ) ^ P0[13];
  assign S[14] = ( G5[13] | ( P5[13] & Cin ) ) ^ P0[14];
  assign S[15] = ( G5[14] | ( P5[14] & Cin ) ) ^ P0[15];
  assign S[16] = ( G5[15] | ( P5[15] & Cin ) ) ^ P0[16];
  assign S[17] = ( G5[16] | ( P5[16] & Cin ) ) ^ P0[17];
  assign S[18] = ( G5[17] | ( P5[17] & Cin ) ) ^ P0[18];
  assign S[19] = ( G5[18] | ( P5[18] & Cin ) ) ^ P0[19];
  assign S[20] = ( G5[19] | ( P5[19] & Cin ) ) ^ P0[20];
  assign S[21] = ( G5[20] | ( P5[20] & Cin ) ) ^ P0[21];
  assign S[22] = ( G5[21] | ( P5[21] & Cin ) ) ^ P0[22];
  assign S[23] = ( G5[22] | ( P5[22] & Cin ) ) ^ P0[23];
  assign S[24] = ( G5[23] | ( P5[23] & Cin ) ) ^ P0[24];
  assign S[25] = ( G5[24] | ( P5[24] & Cin ) ) ^ P0[25];
  assign S[26] = ( G5[25] | ( P5[25] & Cin ) ) ^ P0[26];
  assign S[27] = ( G5[26] | ( P5[26] & Cin ) ) ^ P0[27];
  assign S[28] = G5[27] | ( P5[27] & Cin );
  GPGenerator U0 (G0[1], P0[1], X[1], Y[1]);
  GPGenerator U1 (G0[2], P0[2], X[2], Y[2]);
  GPGenerator U2 (G0[3], P0[3], X[3], Y[3]);
  GPGenerator U3 (G0[4], P0[4], X[4], Y[4]);
  GPGenerator U4 (G0[5], P0[5], X[5], Y[5]);
  GPGenerator U5 (G0[6], P0[6], X[6], Y[6]);
  GPGenerator U6 (G0[7], P0[7], X[7], Y[7]);
  GPGenerator U7 (G0[8], P0[8], X[8], Y[8]);
  GPGenerator U8 (G0[9], P0[9], X[9], Y[9]);
  GPGenerator U9 (G0[10], P0[10], X[10], Y[10]);
  GPGenerator U10 (G0[11], P0[11], X[11], Y[11]);
  GPGenerator U11 (G0[12], P0[12], X[12], Y[12]);
  GPGenerator U12 (G0[13], P0[13], X[13], Y[13]);
  GPGenerator U13 (G0[14], P0[14], X[14], Y[14]);
  GPGenerator U14 (G0[15], P0[15], X[15], Y[15]);
  GPGenerator U15 (G0[16], P0[16], X[16], Y[16]);
  GPGenerator U16 (G0[17], P0[17], X[17], Y[17]);
  GPGenerator U17 (G0[18], P0[18], X[18], Y[18]);
  GPGenerator U18 (G0[19], P0[19], X[19], Y[19]);
  GPGenerator U19 (G0[20], P0[20], X[20], Y[20]);
  GPGenerator U20 (G0[21], P0[21], X[21], Y[21]);
  GPGenerator U21 (G0[22], P0[22], X[22], Y[22]);
  GPGenerator U22 (G0[23], P0[23], X[23], Y[23]);
  GPGenerator U23 (G0[24], P0[24], X[24], Y[24]);
  GPGenerator U24 (G0[25], P0[25], X[25], Y[25]);
  GPGenerator U25 (G0[26], P0[26], X[26], Y[26]);
  GPGenerator U26 (G0[27], P0[27], X[27], Y[27]);
  CarryOperator U27 (G1[2], P1[2], G0[2], P0[2], G0[1], P0[1]);
  CarryOperator U28 (G1[3], P1[3], G0[3], P0[3], G0[2], P0[2]);
  CarryOperator U29 (G1[4], P1[4], G0[4], P0[4], G0[3], P0[3]);
  CarryOperator U30 (G1[5], P1[5], G0[5], P0[5], G0[4], P0[4]);
  CarryOperator U31 (G1[6], P1[6], G0[6], P0[6], G0[5], P0[5]);
  CarryOperator U32 (G1[7], P1[7], G0[7], P0[7], G0[6], P0[6]);
  CarryOperator U33 (G1[8], P1[8], G0[8], P0[8], G0[7], P0[7]);
  CarryOperator U34 (G1[9], P1[9], G0[9], P0[9], G0[8], P0[8]);
  CarryOperator U35 (G1[10], P1[10], G0[10], P0[10], G0[9], P0[9]);
  CarryOperator U36 (G1[11], P1[11], G0[11], P0[11], G0[10], P0[10]);
  CarryOperator U37 (G1[12], P1[12], G0[12], P0[12], G0[11], P0[11]);
  CarryOperator U38 (G1[13], P1[13], G0[13], P0[13], G0[12], P0[12]);
  CarryOperator U39 (G1[14], P1[14], G0[14], P0[14], G0[13], P0[13]);
  CarryOperator U40 (G1[15], P1[15], G0[15], P0[15], G0[14], P0[14]);
  CarryOperator U41 (G1[16], P1[16], G0[16], P0[16], G0[15], P0[15]);
  CarryOperator U42 (G1[17], P1[17], G0[17], P0[17], G0[16], P0[16]);
  CarryOperator U43 (G1[18], P1[18], G0[18], P0[18], G0[17], P0[17]);
  CarryOperator U44 (G1[19], P1[19], G0[19], P0[19], G0[18], P0[18]);
  CarryOperator U45 (G1[20], P1[20], G0[20], P0[20], G0[19], P0[19]);
  CarryOperator U46 (G1[21], P1[21], G0[21], P0[21], G0[20], P0[20]);
  CarryOperator U47 (G1[22], P1[22], G0[22], P0[22], G0[21], P0[21]);
  CarryOperator U48 (G1[23], P1[23], G0[23], P0[23], G0[22], P0[22]);
  CarryOperator U49 (G1[24], P1[24], G0[24], P0[24], G0[23], P0[23]);
  CarryOperator U50 (G1[25], P1[25], G0[25], P0[25], G0[24], P0[24]);
  CarryOperator U51 (G1[26], P1[26], G0[26], P0[26], G0[25], P0[25]);
  CarryOperator U52 (G1[27], P1[27], G0[27], P0[27], G0[26], P0[26]);
  CarryOperator U53 (G2[3], P2[3], G1[3], P1[3], G1[1], P1[1]);
  CarryOperator U54 (G2[4], P2[4], G1[4], P1[4], G1[2], P1[2]);
  CarryOperator U55 (G2[5], P2[5], G1[5], P1[5], G1[3], P1[3]);
  CarryOperator U56 (G2[6], P2[6], G1[6], P1[6], G1[4], P1[4]);
  CarryOperator U57 (G2[7], P2[7], G1[7], P1[7], G1[5], P1[5]);
  CarryOperator U58 (G2[8], P2[8], G1[8], P1[8], G1[6], P1[6]);
  CarryOperator U59 (G2[9], P2[9], G1[9], P1[9], G1[7], P1[7]);
  CarryOperator U60 (G2[10], P2[10], G1[10], P1[10], G1[8], P1[8]);
  CarryOperator U61 (G2[11], P2[11], G1[11], P1[11], G1[9], P1[9]);
  CarryOperator U62 (G2[12], P2[12], G1[12], P1[12], G1[10], P1[10]);
  CarryOperator U63 (G2[13], P2[13], G1[13], P1[13], G1[11], P1[11]);
  CarryOperator U64 (G2[14], P2[14], G1[14], P1[14], G1[12], P1[12]);
  CarryOperator U65 (G2[15], P2[15], G1[15], P1[15], G1[13], P1[13]);
  CarryOperator U66 (G2[16], P2[16], G1[16], P1[16], G1[14], P1[14]);
  CarryOperator U67 (G2[17], P2[17], G1[17], P1[17], G1[15], P1[15]);
  CarryOperator U68 (G2[18], P2[18], G1[18], P1[18], G1[16], P1[16]);
  CarryOperator U69 (G2[19], P2[19], G1[19], P1[19], G1[17], P1[17]);
  CarryOperator U70 (G2[20], P2[20], G1[20], P1[20], G1[18], P1[18]);
  CarryOperator U71 (G2[21], P2[21], G1[21], P1[21], G1[19], P1[19]);
  CarryOperator U72 (G2[22], P2[22], G1[22], P1[22], G1[20], P1[20]);
  CarryOperator U73 (G2[23], P2[23], G1[23], P1[23], G1[21], P1[21]);
  CarryOperator U74 (G2[24], P2[24], G1[24], P1[24], G1[22], P1[22]);
  CarryOperator U75 (G2[25], P2[25], G1[25], P1[25], G1[23], P1[23]);
  CarryOperator U76 (G2[26], P2[26], G1[26], P1[26], G1[24], P1[24]);
  CarryOperator U77 (G2[27], P2[27], G1[27], P1[27], G1[25], P1[25]);
  CarryOperator U78 (G3[5], P3[5], G2[5], P2[5], G2[1], P2[1]);
  CarryOperator U79 (G3[6], P3[6], G2[6], P2[6], G2[2], P2[2]);
  CarryOperator U80 (G3[7], P3[7], G2[7], P2[7], G2[3], P2[3]);
  CarryOperator U81 (G3[8], P3[8], G2[8], P2[8], G2[4], P2[4]);
  CarryOperator U82 (G3[9], P3[9], G2[9], P2[9], G2[5], P2[5]);
  CarryOperator U83 (G3[10], P3[10], G2[10], P2[10], G2[6], P2[6]);
  CarryOperator U84 (G3[11], P3[11], G2[11], P2[11], G2[7], P2[7]);
  CarryOperator U85 (G3[12], P3[12], G2[12], P2[12], G2[8], P2[8]);
  CarryOperator U86 (G3[13], P3[13], G2[13], P2[13], G2[9], P2[9]);
  CarryOperator U87 (G3[14], P3[14], G2[14], P2[14], G2[10], P2[10]);
  CarryOperator U88 (G3[15], P3[15], G2[15], P2[15], G2[11], P2[11]);
  CarryOperator U89 (G3[16], P3[16], G2[16], P2[16], G2[12], P2[12]);
  CarryOperator U90 (G3[17], P3[17], G2[17], P2[17], G2[13], P2[13]);
  CarryOperator U91 (G3[18], P3[18], G2[18], P2[18], G2[14], P2[14]);
  CarryOperator U92 (G3[19], P3[19], G2[19], P2[19], G2[15], P2[15]);
  CarryOperator U93 (G3[20], P3[20], G2[20], P2[20], G2[16], P2[16]);
  CarryOperator U94 (G3[21], P3[21], G2[21], P2[21], G2[17], P2[17]);
  CarryOperator U95 (G3[22], P3[22], G2[22], P2[22], G2[18], P2[18]);
  CarryOperator U96 (G3[23], P3[23], G2[23], P2[23], G2[19], P2[19]);
  CarryOperator U97 (G3[24], P3[24], G2[24], P2[24], G2[20], P2[20]);
  CarryOperator U98 (G3[25], P3[25], G2[25], P2[25], G2[21], P2[21]);
  CarryOperator U99 (G3[26], P3[26], G2[26], P2[26], G2[22], P2[22]);
  CarryOperator U100 (G3[27], P3[27], G2[27], P2[27], G2[23], P2[23]);
  CarryOperator U101 (G4[9], P4[9], G3[9], P3[9], G3[1], P3[1]);
  CarryOperator U102 (G4[10], P4[10], G3[10], P3[10], G3[2], P3[2]);
  CarryOperator U103 (G4[11], P4[11], G3[11], P3[11], G3[3], P3[3]);
  CarryOperator U104 (G4[12], P4[12], G3[12], P3[12], G3[4], P3[4]);
  CarryOperator U105 (G4[13], P4[13], G3[13], P3[13], G3[5], P3[5]);
  CarryOperator U106 (G4[14], P4[14], G3[14], P3[14], G3[6], P3[6]);
  CarryOperator U107 (G4[15], P4[15], G3[15], P3[15], G3[7], P3[7]);
  CarryOperator U108 (G4[16], P4[16], G3[16], P3[16], G3[8], P3[8]);
  CarryOperator U109 (G4[17], P4[17], G3[17], P3[17], G3[9], P3[9]);
  CarryOperator U110 (G4[18], P4[18], G3[18], P3[18], G3[10], P3[10]);
  CarryOperator U111 (G4[19], P4[19], G3[19], P3[19], G3[11], P3[11]);
  CarryOperator U112 (G4[20], P4[20], G3[20], P3[20], G3[12], P3[12]);
  CarryOperator U113 (G4[21], P4[21], G3[21], P3[21], G3[13], P3[13]);
  CarryOperator U114 (G4[22], P4[22], G3[22], P3[22], G3[14], P3[14]);
  CarryOperator U115 (G4[23], P4[23], G3[23], P3[23], G3[15], P3[15]);
  CarryOperator U116 (G4[24], P4[24], G3[24], P3[24], G3[16], P3[16]);
  CarryOperator U117 (G4[25], P4[25], G3[25], P3[25], G3[17], P3[17]);
  CarryOperator U118 (G4[26], P4[26], G3[26], P3[26], G3[18], P3[18]);
  CarryOperator U119 (G4[27], P4[27], G3[27], P3[27], G3[19], P3[19]);
  CarryOperator U120 (G5[17], P5[17], G4[17], P4[17], G4[1], P4[1]);
  CarryOperator U121 (G5[18], P5[18], G4[18], P4[18], G4[2], P4[2]);
  CarryOperator U122 (G5[19], P5[19], G4[19], P4[19], G4[3], P4[3]);
  CarryOperator U123 (G5[20], P5[20], G4[20], P4[20], G4[4], P4[4]);
  CarryOperator U124 (G5[21], P5[21], G4[21], P4[21], G4[5], P4[5]);
  CarryOperator U125 (G5[22], P5[22], G4[22], P4[22], G4[6], P4[6]);
  CarryOperator U126 (G5[23], P5[23], G4[23], P4[23], G4[7], P4[7]);
  CarryOperator U127 (G5[24], P5[24], G4[24], P4[24], G4[8], P4[8]);
  CarryOperator U128 (G5[25], P5[25], G4[25], P4[25], G4[9], P4[9]);
  CarryOperator U129 (G5[26], P5[26], G4[26], P4[26], G4[10], P4[10]);
  CarryOperator U130 (G5[27], P5[27], G4[27], P4[27], G4[11], P4[11]);
endmodule

module UBZero_1_1(O);
  output [1:1] O;
  assign O[1] = 0;
endmodule

module Multiplier_13_0_1000(P, IN1, IN2);
  output [27:0] P;
  input [13:0] IN1;
  input [13:0] IN2;
  wire [28:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  assign P[12] = W[12];
  assign P[13] = W[13];
  assign P[14] = W[14];
  assign P[15] = W[15];
  assign P[16] = W[16];
  assign P[17] = W[17];
  assign P[18] = W[18];
  assign P[19] = W[19];
  assign P[20] = W[20];
  assign P[21] = W[21];
  assign P[22] = W[22];
  assign P[23] = W[23];
  assign P[24] = W[24];
  assign P[25] = W[25];
  assign P[26] = W[26];
  assign P[27] = W[27];
  MultUB_STD_D73_KS000 U0 (W, IN1, IN2);
endmodule

module D7_3CTR_13_0_14_1000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13);
  output [27:0] S1;
  output [26:1] S2;
  input [13:0] PP0;
  input [14:1] PP1;
  input [23:10] PP10;
  input [24:11] PP11;
  input [25:12] PP12;
  input [26:13] PP13;
  input [15:2] PP2;
  input [16:3] PP3;
  input [17:4] PP4;
  input [18:5] PP5;
  input [19:6] PP6;
  input [20:7] PP7;
  input [21:8] PP8;
  input [22:9] PP9;
  wire [26:0] W0;
  wire [25:1] W1;
  wire [24:2] W2;
  wire [23:3] W3;
  wire [22:4] W4;
  wire [22:5] W5;
  wire [21:6] W6;
  UBHA_7 U0 (W5[8], W6[7], PP0[7], PP1[7]);
  UB4_3C8 U1 (W4[10], W5[9], W6[8], PP0[8], PP1[8], PP2[8], PP3[8]);
  UB5_3C9 U2 (W3[11], W5[10], W6[9], PP0[9], PP1[9], PP2[9], PP3[9], PP4[9]);
  UB7_3C10 U3 (W2[12], W4[11], W6[10], PP0[10], PP1[10], PP2[10], PP3[10], PP4[10], PP5[10], PP6[10]);
  UB7_3C11 U4 (W2[13], W3[12], W5[11], PP0[11], PP1[11], PP2[11], PP3[11], PP4[11], PP5[11], PP6[11]);
  UBHA_11 U5 (W4[12], W6[11], PP7[11], PP8[11]);
  UB7_3C12 U6 (W1[14], W3[13], W5[12], PP0[12], PP1[12], PP2[12], PP3[12], PP4[12], PP5[12], PP6[12]);
  UB4_3C12 U7 (W2[14], W4[13], W6[12], PP7[12], PP8[12], PP9[12], PP10[12]);
  UB7_3C13 U8 (W1[15], W3[14], W5[13], PP0[13], PP1[13], PP2[13], PP3[13], PP4[13], PP5[13], PP6[13]);
  UB5_3C13 U9 (W2[15], W4[14], W6[13], PP7[13], PP8[13], PP9[13], PP10[13], PP11[13]);
  UB7_3C14 U10 (W1[16], W3[15], W5[14], PP1[14], PP2[14], PP3[14], PP4[14], PP5[14], PP6[14], PP7[14]);
  UB5_3C14 U11 (W2[16], W4[15], W6[14], PP8[14], PP9[14], PP10[14], PP11[14], PP12[14]);
  UB7_3C15 U12 (W1[17], W3[16], W5[15], PP2[15], PP3[15], PP4[15], PP5[15], PP6[15], PP7[15], PP8[15]);
  UB4_3C15 U13 (W2[17], W4[16], W6[15], PP9[15], PP10[15], PP11[15], PP12[15]);
  UB7_3C16 U14 (W3[18], W3[17], W5[16], PP3[16], PP4[16], PP5[16], PP6[16], PP7[16], PP8[16], PP9[16]);
  UBFA_16 U15 (W4[17], W6[16], PP10[16], PP11[16], PP12[16]);
  UB7_3C17 U16 (W4[19], W4[18], W5[17], PP4[17], PP5[17], PP6[17], PP7[17], PP8[17], PP9[17], PP10[17]);
  UBHA_17 U17 (W5[18], W6[17], PP11[17], PP12[17]);
  UB6_3C18 U18 (W4[20], W5[19], W6[18], PP5[18], PP6[18], PP7[18], PP8[18], PP9[18], PP10[18]);
  UB4_3C19 U19 (W4[21], W5[20], W6[19], PP6[19], PP7[19], PP8[19], PP9[19]);
  UBFA_20 U20 (W5[21], W6[20], PP7[20], PP8[20], PP9[20]);
  UBHA_21 U21 (W5[22], W6[21], PP8[21], PP9[21]);
  UBCON_6_0 U22 (W0[6:0], PP0[6:0]);
  UB1DCON_7 U23 (W0[7], PP2[7]);
  UB1DCON_8 U24 (W0[8], PP4[8]);
  UB1DCON_9 U25 (W0[9], PP5[9]);
  UB1DCON_10 U26 (W0[10], PP7[10]);
  UB1DCON_11 U27 (W0[11], PP9[11]);
  UB1DCON_12 U28 (W0[12], PP11[12]);
  UB1DCON_13 U29 (W0[13], PP12[13]);
  UBCON_17_14 U30 (W0[17:14], PP13[17:14]);
  UB1DCON_18 U31 (W0[18], PP11[18]);
  UBCON_21_19 U32 (W0[21:19], PP10[21:19]);
  UB1DCON_22 U33 (W0[22], PP9[22]);
  UB1DCON_23 U34 (W0[23], PP10[23]);
  UB1DCON_24 U35 (W0[24], PP11[24]);
  UB1DCON_25 U36 (W0[25], PP12[25]);
  UB1DCON_26 U37 (W0[26], PP13[26]);
  UBCON_6_1 U38 (W1[6:1], PP1[6:1]);
  UB1DCON_7 U39 (W1[7], PP3[7]);
  UB1DCON_8 U40 (W1[8], PP5[8]);
  UB1DCON_9 U41 (W1[9], PP6[9]);
  UB1DCON_10 U42 (W1[10], PP8[10]);
  UB1DCON_11 U43 (W1[11], PP10[11]);
  UB1DCON_12 U44 (W1[12], PP12[12]);
  UB1DCON_13 U45 (W1[13], PP13[13]);
  UB1DCON_18 U46 (W1[18], PP12[18]);
  UBCON_21_19 U47 (W1[21:19], PP11[21:19]);
  UB1DCON_22 U48 (W1[22], PP10[22]);
  UB1DCON_23 U49 (W1[23], PP11[23]);
  UB1DCON_24 U50 (W1[24], PP12[24]);
  UB1DCON_25 U51 (W1[25], PP13[25]);
  UBCON_6_2 U52 (W2[6:2], PP2[6:2]);
  UB1DCON_7 U53 (W2[7], PP4[7]);
  UB1DCON_8 U54 (W2[8], PP6[8]);
  UB1DCON_9 U55 (W2[9], PP7[9]);
  UB1DCON_10 U56 (W2[10], PP9[10]);
  UB1DCON_11 U57 (W2[11], PP11[11]);
  UB1DCON_18 U58 (W2[18], PP13[18]);
  UBCON_21_19 U59 (W2[21:19], PP12[21:19]);
  UB1DCON_22 U60 (W2[22], PP11[22]);
  UB1DCON_23 U61 (W2[23], PP12[23]);
  UB1DCON_24 U62 (W2[24], PP13[24]);
  UBCON_6_3 U63 (W3[6:3], PP3[6:3]);
  UB1DCON_7 U64 (W3[7], PP5[7]);
  UB1DCON_8 U65 (W3[8], PP7[8]);
  UB1DCON_9 U66 (W3[9], PP8[9]);
  UB1DCON_10 U67 (W3[10], PP10[10]);
  UBCON_21_19 U68 (W3[21:19], PP13[21:19]);
  UB1DCON_22 U69 (W3[22], PP12[22]);
  UB1DCON_23 U70 (W3[23], PP13[23]);
  UBCON_6_4 U71 (W4[6:4], PP4[6:4]);
  UB1DCON_7 U72 (W4[7], PP6[7]);
  UB1DCON_8 U73 (W4[8], PP8[8]);
  UB1DCON_9 U74 (W4[9], PP9[9]);
  UB1DCON_22 U75 (W4[22], PP13[22]);
  UBCON_6_5 U76 (W5[6:5], PP5[6:5]);
  UB1DCON_7 U77 (W5[7], PP7[7]);
  UB1DCON_6 U78 (W6[6], PP6[6]);
  D7_3CTR_26_0_25_1000 U79 (S1, S2, W0, W1, W2, W3, W4, W5, W6);
endmodule

module D7_3CTR_26_0_25_1000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6);
  output [27:0] S1;
  output [26:1] S2;
  input [26:0] PP0;
  input [25:1] PP1;
  input [24:2] PP2;
  input [23:3] PP3;
  input [22:4] PP4;
  input [22:5] PP5;
  input [21:6] PP6;
  wire [26:0] W0;
  wire [26:1] W1;
  wire [25:2] W2;
  UBHA_3 U0 (W1[4], W2[3], PP0[3], PP1[3]);
  UB4_3C4 U1 (W0[6], W1[5], W2[4], PP0[4], PP1[4], PP2[4], PP3[4]);
  UB5_3C5 U2 (W0[7], W1[6], W2[5], PP0[5], PP1[5], PP2[5], PP3[5], PP4[5]);
  UB7_3C6 U3 (W0[8], W1[7], W2[6], PP0[6], PP1[6], PP2[6], PP3[6], PP4[6], PP5[6], PP6[6]);
  UB7_3C7 U4 (W0[9], W1[8], W2[7], PP0[7], PP1[7], PP2[7], PP3[7], PP4[7], PP5[7], PP6[7]);
  UB7_3C8 U5 (W0[10], W1[9], W2[8], PP0[8], PP1[8], PP2[8], PP3[8], PP4[8], PP5[8], PP6[8]);
  UB7_3C9 U6 (W0[11], W1[10], W2[9], PP0[9], PP1[9], PP2[9], PP3[9], PP4[9], PP5[9], PP6[9]);
  UB7_3C10 U7 (W0[12], W1[11], W2[10], PP0[10], PP1[10], PP2[10], PP3[10], PP4[10], PP5[10], PP6[10]);
  UB7_3C11 U8 (W0[13], W1[12], W2[11], PP0[11], PP1[11], PP2[11], PP3[11], PP4[11], PP5[11], PP6[11]);
  UB7_3C12 U9 (W0[14], W1[13], W2[12], PP0[12], PP1[12], PP2[12], PP3[12], PP4[12], PP5[12], PP6[12]);
  UB7_3C13 U10 (W0[15], W1[14], W2[13], PP0[13], PP1[13], PP2[13], PP3[13], PP4[13], PP5[13], PP6[13]);
  UB7_3C14 U11 (W0[16], W1[15], W2[14], PP0[14], PP1[14], PP2[14], PP3[14], PP4[14], PP5[14], PP6[14]);
  UB7_3C15 U12 (W0[17], W1[16], W2[15], PP0[15], PP1[15], PP2[15], PP3[15], PP4[15], PP5[15], PP6[15]);
  UB7_3C16 U13 (W0[18], W1[17], W2[16], PP0[16], PP1[16], PP2[16], PP3[16], PP4[16], PP5[16], PP6[16]);
  UB7_3C17 U14 (W0[19], W1[18], W2[17], PP0[17], PP1[17], PP2[17], PP3[17], PP4[17], PP5[17], PP6[17]);
  UB7_3C18 U15 (W0[20], W1[19], W2[18], PP0[18], PP1[18], PP2[18], PP3[18], PP4[18], PP5[18], PP6[18]);
  UB7_3C19 U16 (W0[21], W1[20], W2[19], PP0[19], PP1[19], PP2[19], PP3[19], PP4[19], PP5[19], PP6[19]);
  UB7_3C20 U17 (W0[22], W1[21], W2[20], PP0[20], PP1[20], PP2[20], PP3[20], PP4[20], PP5[20], PP6[20]);
  UB7_3C21 U18 (W0[23], W1[22], W2[21], PP0[21], PP1[21], PP2[21], PP3[21], PP4[21], PP5[21], PP6[21]);
  UB6_3C22 U19 (W0[24], W1[23], W2[22], PP0[22], PP1[22], PP2[22], PP3[22], PP4[22], PP5[22]);
  UB4_3C23 U20 (W0[25], W1[24], W2[23], PP0[23], PP1[23], PP2[23], PP3[23]);
  UBFA_24 U21 (W1[25], W2[24], PP0[24], PP1[24], PP2[24]);
  UBHA_25 U22 (W1[26], W2[25], PP0[25], PP1[25]);
  UBCON_2_0 U23 (W0[2:0], PP0[2:0]);
  UB1DCON_3 U24 (W0[3], PP2[3]);
  UB1DCON_4 U25 (W0[4], PP4[4]);
  UB1DCON_5 U26 (W0[5], PP5[5]);
  UB1DCON_26 U27 (W0[26], PP0[26]);
  UBCON_2_1 U28 (W1[2:1], PP1[2:1]);
  UB1DCON_3 U29 (W1[3], PP3[3]);
  UB1DCON_2 U30 (W2[2], PP2[2]);
  D7_3CTR_26_0_26_1000 U31 (S1, S2, W0, W1, W2);
endmodule

module D7_3CTR_26_0_26_1000 (S1, S2, PP0, PP1, PP2);
  output [27:0] S1;
  output [26:1] S2;
  input [26:0] PP0;
  input [26:1] PP1;
  input [25:2] PP2;
  wire [27:0] W0;
  wire [26:1] W1;
  UBHA_2 U0 (W0[3], W1[2], PP0[2], PP1[2]);
  UBFA_3 U1 (W0[4], W1[3], PP0[3], PP1[3], PP2[3]);
  UBFA_4 U2 (W0[5], W1[4], PP0[4], PP1[4], PP2[4]);
  UBFA_5 U3 (W0[6], W1[5], PP0[5], PP1[5], PP2[5]);
  UBFA_6 U4 (W0[7], W1[6], PP0[6], PP1[6], PP2[6]);
  UBFA_7 U5 (W0[8], W1[7], PP0[7], PP1[7], PP2[7]);
  UBFA_8 U6 (W0[9], W1[8], PP0[8], PP1[8], PP2[8]);
  UBFA_9 U7 (W0[10], W1[9], PP0[9], PP1[9], PP2[9]);
  UBFA_10 U8 (W0[11], W1[10], PP0[10], PP1[10], PP2[10]);
  UBFA_11 U9 (W0[12], W1[11], PP0[11], PP1[11], PP2[11]);
  UBFA_12 U10 (W0[13], W1[12], PP0[12], PP1[12], PP2[12]);
  UBFA_13 U11 (W0[14], W1[13], PP0[13], PP1[13], PP2[13]);
  UBFA_14 U12 (W0[15], W1[14], PP0[14], PP1[14], PP2[14]);
  UBFA_15 U13 (W0[16], W1[15], PP0[15], PP1[15], PP2[15]);
  UBFA_16 U14 (W0[17], W1[16], PP0[16], PP1[16], PP2[16]);
  UBFA_17 U15 (W0[18], W1[17], PP0[17], PP1[17], PP2[17]);
  UBFA_18 U16 (W0[19], W1[18], PP0[18], PP1[18], PP2[18]);
  UBFA_19 U17 (W0[20], W1[19], PP0[19], PP1[19], PP2[19]);
  UBFA_20 U18 (W0[21], W1[20], PP0[20], PP1[20], PP2[20]);
  UBFA_21 U19 (W0[22], W1[21], PP0[21], PP1[21], PP2[21]);
  UBFA_22 U20 (W0[23], W1[22], PP0[22], PP1[22], PP2[22]);
  UBFA_23 U21 (W0[24], W1[23], PP0[23], PP1[23], PP2[23]);
  UBFA_24 U22 (W0[25], W1[24], PP0[24], PP1[24], PP2[24]);
  UBFA_25 U23 (W0[26], W1[25], PP0[25], PP1[25], PP2[25]);
  UBHA_26 U24 (W0[27], W1[26], PP0[26], PP1[26]);
  UBCON_1_0 U25 (W0[1:0], PP0[1:0]);
  UB1DCON_2 U26 (W0[2], PP2[2]);
  UB1DCON_1 U27 (W1[1], PP1[1]);
  D7_3CTR_27_0_26_1 U28 (S1, S2, W0, W1);
endmodule

module D7_3CTR_27_0_26_1 (S1, S2, PP0, PP1);
  output [27:0] S1;
  output [26:1] S2;
  input [27:0] PP0;
  input [26:1] PP1;
  UBCON_27_0 U0 (S1, PP0);
  UBCON_26_1 U1 (S2, PP1);
endmodule

module MultUB_STD_D73_KS000 (P, IN1, IN2);
  output [28:0] P;
  input [13:0] IN1;
  input [13:0] IN2;
  wire [13:0] PP0;
  wire [14:1] PP1;
  wire [23:10] PP10;
  wire [24:11] PP11;
  wire [25:12] PP12;
  wire [26:13] PP13;
  wire [15:2] PP2;
  wire [16:3] PP3;
  wire [17:4] PP4;
  wire [18:5] PP5;
  wire [19:6] PP6;
  wire [20:7] PP7;
  wire [21:8] PP8;
  wire [22:9] PP9;
  wire [27:0] S1;
  wire [26:1] S2;
  UBPPG_13_0_13_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, IN1, IN2);
  D7_3CTR_13_0_14_1000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13);
  UBKSA_27_0_26_1 U2 (P, S1, S2);
endmodule

module UBCON_17_14 (O, I);
  output [17:14] O;
  input [17:14] I;
  UB1DCON_14 U0 (O[14], I[14]);
  UB1DCON_15 U1 (O[15], I[15]);
  UB1DCON_16 U2 (O[16], I[16]);
  UB1DCON_17 U3 (O[17], I[17]);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_21_19 (O, I);
  output [21:19] O;
  input [21:19] I;
  UB1DCON_19 U0 (O[19], I[19]);
  UB1DCON_20 U1 (O[20], I[20]);
  UB1DCON_21 U2 (O[21], I[21]);
endmodule

module UBCON_26_1 (O, I);
  output [26:1] O;
  input [26:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
  UB1DCON_6 U5 (O[6], I[6]);
  UB1DCON_7 U6 (O[7], I[7]);
  UB1DCON_8 U7 (O[8], I[8]);
  UB1DCON_9 U8 (O[9], I[9]);
  UB1DCON_10 U9 (O[10], I[10]);
  UB1DCON_11 U10 (O[11], I[11]);
  UB1DCON_12 U11 (O[12], I[12]);
  UB1DCON_13 U12 (O[13], I[13]);
  UB1DCON_14 U13 (O[14], I[14]);
  UB1DCON_15 U14 (O[15], I[15]);
  UB1DCON_16 U15 (O[16], I[16]);
  UB1DCON_17 U16 (O[17], I[17]);
  UB1DCON_18 U17 (O[18], I[18]);
  UB1DCON_19 U18 (O[19], I[19]);
  UB1DCON_20 U19 (O[20], I[20]);
  UB1DCON_21 U20 (O[21], I[21]);
  UB1DCON_22 U21 (O[22], I[22]);
  UB1DCON_23 U22 (O[23], I[23]);
  UB1DCON_24 U23 (O[24], I[24]);
  UB1DCON_25 U24 (O[25], I[25]);
  UB1DCON_26 U25 (O[26], I[26]);
endmodule

module UBCON_27_0 (O, I);
  output [27:0] O;
  input [27:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
  UB1DCON_13 U13 (O[13], I[13]);
  UB1DCON_14 U14 (O[14], I[14]);
  UB1DCON_15 U15 (O[15], I[15]);
  UB1DCON_16 U16 (O[16], I[16]);
  UB1DCON_17 U17 (O[17], I[17]);
  UB1DCON_18 U18 (O[18], I[18]);
  UB1DCON_19 U19 (O[19], I[19]);
  UB1DCON_20 U20 (O[20], I[20]);
  UB1DCON_21 U21 (O[21], I[21]);
  UB1DCON_22 U22 (O[22], I[22]);
  UB1DCON_23 U23 (O[23], I[23]);
  UB1DCON_24 U24 (O[24], I[24]);
  UB1DCON_25 U25 (O[25], I[25]);
  UB1DCON_26 U26 (O[26], I[26]);
  UB1DCON_27 U27 (O[27], I[27]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBCON_2_1 (O, I);
  output [2:1] O;
  input [2:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
endmodule

module UBCON_6_0 (O, I);
  output [6:0] O;
  input [6:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
endmodule

module UBCON_6_1 (O, I);
  output [6:1] O;
  input [6:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
  UB1DCON_6 U5 (O[6], I[6]);
endmodule

module UBCON_6_2 (O, I);
  output [6:2] O;
  input [6:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
  UB1DCON_6 U4 (O[6], I[6]);
endmodule

module UBCON_6_3 (O, I);
  output [6:3] O;
  input [6:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
  UB1DCON_6 U3 (O[6], I[6]);
endmodule

module UBCON_6_4 (O, I);
  output [6:4] O;
  input [6:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
endmodule

module UBCON_6_5 (O, I);
  output [6:5] O;
  input [6:5] I;
  UB1DCON_5 U0 (O[5], I[5]);
  UB1DCON_6 U1 (O[6], I[6]);
endmodule

module UBExtender_26_1_2000 (O, I);
  output [27:1] O;
  input [26:1] I;
  UBCON_26_1 U0 (O[26:1], I[26:1]);
  UBZero_27_27 U1 (O[27]);
endmodule

module UBKSA_27_0_26_1 (S, X, Y);
  output [28:0] S;
  input [27:0] X;
  input [26:1] Y;
  wire [27:1] Z;
  UBExtender_26_1_2000 U0 (Z[27:1], Y[26:1]);
  UBPureKSA_27_1 U1 (S[28:1], X[27:1], Z[27:1]);
  UB1DCON_0 U2 (S[0], X[0]);
endmodule

module UBPPG_13_0_13_0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, IN1, IN2);
  output [13:0] PP0;
  output [14:1] PP1;
  output [23:10] PP10;
  output [24:11] PP11;
  output [25:12] PP12;
  output [26:13] PP13;
  output [15:2] PP2;
  output [16:3] PP3;
  output [17:4] PP4;
  output [18:5] PP5;
  output [19:6] PP6;
  output [20:7] PP7;
  output [21:8] PP8;
  output [22:9] PP9;
  input [13:0] IN1;
  input [13:0] IN2;
  UBVPPG_13_0_0 U0 (PP0, IN1, IN2[0]);
  UBVPPG_13_0_1 U1 (PP1, IN1, IN2[1]);
  UBVPPG_13_0_2 U2 (PP2, IN1, IN2[2]);
  UBVPPG_13_0_3 U3 (PP3, IN1, IN2[3]);
  UBVPPG_13_0_4 U4 (PP4, IN1, IN2[4]);
  UBVPPG_13_0_5 U5 (PP5, IN1, IN2[5]);
  UBVPPG_13_0_6 U6 (PP6, IN1, IN2[6]);
  UBVPPG_13_0_7 U7 (PP7, IN1, IN2[7]);
  UBVPPG_13_0_8 U8 (PP8, IN1, IN2[8]);
  UBVPPG_13_0_9 U9 (PP9, IN1, IN2[9]);
  UBVPPG_13_0_10 U10 (PP10, IN1, IN2[10]);
  UBVPPG_13_0_11 U11 (PP11, IN1, IN2[11]);
  UBVPPG_13_0_12 U12 (PP12, IN1, IN2[12]);
  UBVPPG_13_0_13 U13 (PP13, IN1, IN2[13]);
endmodule

module UBPureKSA_27_1 (S, X, Y);
  output [28:1] S;
  input [27:1] X;
  input [27:1] Y;
  wire C;
  UBPriKSA_27_1 U0 (S, X, Y, C);
  UBZero_1_1 U1 (C);
endmodule

module UBVPPG_13_0_0 (O, IN1, IN2);
  output [13:0] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
  UB1BPPG_6_0 U6 (O[6], IN1[6], IN2);
  UB1BPPG_7_0 U7 (O[7], IN1[7], IN2);
  UB1BPPG_8_0 U8 (O[8], IN1[8], IN2);
  UB1BPPG_9_0 U9 (O[9], IN1[9], IN2);
  UB1BPPG_10_0 U10 (O[10], IN1[10], IN2);
  UB1BPPG_11_0 U11 (O[11], IN1[11], IN2);
  UB1BPPG_12_0 U12 (O[12], IN1[12], IN2);
  UB1BPPG_13_0 U13 (O[13], IN1[13], IN2);
endmodule

module UBVPPG_13_0_1 (O, IN1, IN2);
  output [14:1] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_1 U0 (O[1], IN1[0], IN2);
  UB1BPPG_1_1 U1 (O[2], IN1[1], IN2);
  UB1BPPG_2_1 U2 (O[3], IN1[2], IN2);
  UB1BPPG_3_1 U3 (O[4], IN1[3], IN2);
  UB1BPPG_4_1 U4 (O[5], IN1[4], IN2);
  UB1BPPG_5_1 U5 (O[6], IN1[5], IN2);
  UB1BPPG_6_1 U6 (O[7], IN1[6], IN2);
  UB1BPPG_7_1 U7 (O[8], IN1[7], IN2);
  UB1BPPG_8_1 U8 (O[9], IN1[8], IN2);
  UB1BPPG_9_1 U9 (O[10], IN1[9], IN2);
  UB1BPPG_10_1 U10 (O[11], IN1[10], IN2);
  UB1BPPG_11_1 U11 (O[12], IN1[11], IN2);
  UB1BPPG_12_1 U12 (O[13], IN1[12], IN2);
  UB1BPPG_13_1 U13 (O[14], IN1[13], IN2);
endmodule

module UBVPPG_13_0_10 (O, IN1, IN2);
  output [23:10] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_10 U0 (O[10], IN1[0], IN2);
  UB1BPPG_1_10 U1 (O[11], IN1[1], IN2);
  UB1BPPG_2_10 U2 (O[12], IN1[2], IN2);
  UB1BPPG_3_10 U3 (O[13], IN1[3], IN2);
  UB1BPPG_4_10 U4 (O[14], IN1[4], IN2);
  UB1BPPG_5_10 U5 (O[15], IN1[5], IN2);
  UB1BPPG_6_10 U6 (O[16], IN1[6], IN2);
  UB1BPPG_7_10 U7 (O[17], IN1[7], IN2);
  UB1BPPG_8_10 U8 (O[18], IN1[8], IN2);
  UB1BPPG_9_10 U9 (O[19], IN1[9], IN2);
  UB1BPPG_10_10 U10 (O[20], IN1[10], IN2);
  UB1BPPG_11_10 U11 (O[21], IN1[11], IN2);
  UB1BPPG_12_10 U12 (O[22], IN1[12], IN2);
  UB1BPPG_13_10 U13 (O[23], IN1[13], IN2);
endmodule

module UBVPPG_13_0_11 (O, IN1, IN2);
  output [24:11] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_11 U0 (O[11], IN1[0], IN2);
  UB1BPPG_1_11 U1 (O[12], IN1[1], IN2);
  UB1BPPG_2_11 U2 (O[13], IN1[2], IN2);
  UB1BPPG_3_11 U3 (O[14], IN1[3], IN2);
  UB1BPPG_4_11 U4 (O[15], IN1[4], IN2);
  UB1BPPG_5_11 U5 (O[16], IN1[5], IN2);
  UB1BPPG_6_11 U6 (O[17], IN1[6], IN2);
  UB1BPPG_7_11 U7 (O[18], IN1[7], IN2);
  UB1BPPG_8_11 U8 (O[19], IN1[8], IN2);
  UB1BPPG_9_11 U9 (O[20], IN1[9], IN2);
  UB1BPPG_10_11 U10 (O[21], IN1[10], IN2);
  UB1BPPG_11_11 U11 (O[22], IN1[11], IN2);
  UB1BPPG_12_11 U12 (O[23], IN1[12], IN2);
  UB1BPPG_13_11 U13 (O[24], IN1[13], IN2);
endmodule

module UBVPPG_13_0_12 (O, IN1, IN2);
  output [25:12] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_12 U0 (O[12], IN1[0], IN2);
  UB1BPPG_1_12 U1 (O[13], IN1[1], IN2);
  UB1BPPG_2_12 U2 (O[14], IN1[2], IN2);
  UB1BPPG_3_12 U3 (O[15], IN1[3], IN2);
  UB1BPPG_4_12 U4 (O[16], IN1[4], IN2);
  UB1BPPG_5_12 U5 (O[17], IN1[5], IN2);
  UB1BPPG_6_12 U6 (O[18], IN1[6], IN2);
  UB1BPPG_7_12 U7 (O[19], IN1[7], IN2);
  UB1BPPG_8_12 U8 (O[20], IN1[8], IN2);
  UB1BPPG_9_12 U9 (O[21], IN1[9], IN2);
  UB1BPPG_10_12 U10 (O[22], IN1[10], IN2);
  UB1BPPG_11_12 U11 (O[23], IN1[11], IN2);
  UB1BPPG_12_12 U12 (O[24], IN1[12], IN2);
  UB1BPPG_13_12 U13 (O[25], IN1[13], IN2);
endmodule

module UBVPPG_13_0_13 (O, IN1, IN2);
  output [26:13] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_13 U0 (O[13], IN1[0], IN2);
  UB1BPPG_1_13 U1 (O[14], IN1[1], IN2);
  UB1BPPG_2_13 U2 (O[15], IN1[2], IN2);
  UB1BPPG_3_13 U3 (O[16], IN1[3], IN2);
  UB1BPPG_4_13 U4 (O[17], IN1[4], IN2);
  UB1BPPG_5_13 U5 (O[18], IN1[5], IN2);
  UB1BPPG_6_13 U6 (O[19], IN1[6], IN2);
  UB1BPPG_7_13 U7 (O[20], IN1[7], IN2);
  UB1BPPG_8_13 U8 (O[21], IN1[8], IN2);
  UB1BPPG_9_13 U9 (O[22], IN1[9], IN2);
  UB1BPPG_10_13 U10 (O[23], IN1[10], IN2);
  UB1BPPG_11_13 U11 (O[24], IN1[11], IN2);
  UB1BPPG_12_13 U12 (O[25], IN1[12], IN2);
  UB1BPPG_13_13 U13 (O[26], IN1[13], IN2);
endmodule

module UBVPPG_13_0_2 (O, IN1, IN2);
  output [15:2] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
  UB1BPPG_6_2 U6 (O[8], IN1[6], IN2);
  UB1BPPG_7_2 U7 (O[9], IN1[7], IN2);
  UB1BPPG_8_2 U8 (O[10], IN1[8], IN2);
  UB1BPPG_9_2 U9 (O[11], IN1[9], IN2);
  UB1BPPG_10_2 U10 (O[12], IN1[10], IN2);
  UB1BPPG_11_2 U11 (O[13], IN1[11], IN2);
  UB1BPPG_12_2 U12 (O[14], IN1[12], IN2);
  UB1BPPG_13_2 U13 (O[15], IN1[13], IN2);
endmodule

module UBVPPG_13_0_3 (O, IN1, IN2);
  output [16:3] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_3 U0 (O[3], IN1[0], IN2);
  UB1BPPG_1_3 U1 (O[4], IN1[1], IN2);
  UB1BPPG_2_3 U2 (O[5], IN1[2], IN2);
  UB1BPPG_3_3 U3 (O[6], IN1[3], IN2);
  UB1BPPG_4_3 U4 (O[7], IN1[4], IN2);
  UB1BPPG_5_3 U5 (O[8], IN1[5], IN2);
  UB1BPPG_6_3 U6 (O[9], IN1[6], IN2);
  UB1BPPG_7_3 U7 (O[10], IN1[7], IN2);
  UB1BPPG_8_3 U8 (O[11], IN1[8], IN2);
  UB1BPPG_9_3 U9 (O[12], IN1[9], IN2);
  UB1BPPG_10_3 U10 (O[13], IN1[10], IN2);
  UB1BPPG_11_3 U11 (O[14], IN1[11], IN2);
  UB1BPPG_12_3 U12 (O[15], IN1[12], IN2);
  UB1BPPG_13_3 U13 (O[16], IN1[13], IN2);
endmodule

module UBVPPG_13_0_4 (O, IN1, IN2);
  output [17:4] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
  UB1BPPG_6_4 U6 (O[10], IN1[6], IN2);
  UB1BPPG_7_4 U7 (O[11], IN1[7], IN2);
  UB1BPPG_8_4 U8 (O[12], IN1[8], IN2);
  UB1BPPG_9_4 U9 (O[13], IN1[9], IN2);
  UB1BPPG_10_4 U10 (O[14], IN1[10], IN2);
  UB1BPPG_11_4 U11 (O[15], IN1[11], IN2);
  UB1BPPG_12_4 U12 (O[16], IN1[12], IN2);
  UB1BPPG_13_4 U13 (O[17], IN1[13], IN2);
endmodule

module UBVPPG_13_0_5 (O, IN1, IN2);
  output [18:5] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_5 U0 (O[5], IN1[0], IN2);
  UB1BPPG_1_5 U1 (O[6], IN1[1], IN2);
  UB1BPPG_2_5 U2 (O[7], IN1[2], IN2);
  UB1BPPG_3_5 U3 (O[8], IN1[3], IN2);
  UB1BPPG_4_5 U4 (O[9], IN1[4], IN2);
  UB1BPPG_5_5 U5 (O[10], IN1[5], IN2);
  UB1BPPG_6_5 U6 (O[11], IN1[6], IN2);
  UB1BPPG_7_5 U7 (O[12], IN1[7], IN2);
  UB1BPPG_8_5 U8 (O[13], IN1[8], IN2);
  UB1BPPG_9_5 U9 (O[14], IN1[9], IN2);
  UB1BPPG_10_5 U10 (O[15], IN1[10], IN2);
  UB1BPPG_11_5 U11 (O[16], IN1[11], IN2);
  UB1BPPG_12_5 U12 (O[17], IN1[12], IN2);
  UB1BPPG_13_5 U13 (O[18], IN1[13], IN2);
endmodule

module UBVPPG_13_0_6 (O, IN1, IN2);
  output [19:6] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_6 U0 (O[6], IN1[0], IN2);
  UB1BPPG_1_6 U1 (O[7], IN1[1], IN2);
  UB1BPPG_2_6 U2 (O[8], IN1[2], IN2);
  UB1BPPG_3_6 U3 (O[9], IN1[3], IN2);
  UB1BPPG_4_6 U4 (O[10], IN1[4], IN2);
  UB1BPPG_5_6 U5 (O[11], IN1[5], IN2);
  UB1BPPG_6_6 U6 (O[12], IN1[6], IN2);
  UB1BPPG_7_6 U7 (O[13], IN1[7], IN2);
  UB1BPPG_8_6 U8 (O[14], IN1[8], IN2);
  UB1BPPG_9_6 U9 (O[15], IN1[9], IN2);
  UB1BPPG_10_6 U10 (O[16], IN1[10], IN2);
  UB1BPPG_11_6 U11 (O[17], IN1[11], IN2);
  UB1BPPG_12_6 U12 (O[18], IN1[12], IN2);
  UB1BPPG_13_6 U13 (O[19], IN1[13], IN2);
endmodule

module UBVPPG_13_0_7 (O, IN1, IN2);
  output [20:7] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_7 U0 (O[7], IN1[0], IN2);
  UB1BPPG_1_7 U1 (O[8], IN1[1], IN2);
  UB1BPPG_2_7 U2 (O[9], IN1[2], IN2);
  UB1BPPG_3_7 U3 (O[10], IN1[3], IN2);
  UB1BPPG_4_7 U4 (O[11], IN1[4], IN2);
  UB1BPPG_5_7 U5 (O[12], IN1[5], IN2);
  UB1BPPG_6_7 U6 (O[13], IN1[6], IN2);
  UB1BPPG_7_7 U7 (O[14], IN1[7], IN2);
  UB1BPPG_8_7 U8 (O[15], IN1[8], IN2);
  UB1BPPG_9_7 U9 (O[16], IN1[9], IN2);
  UB1BPPG_10_7 U10 (O[17], IN1[10], IN2);
  UB1BPPG_11_7 U11 (O[18], IN1[11], IN2);
  UB1BPPG_12_7 U12 (O[19], IN1[12], IN2);
  UB1BPPG_13_7 U13 (O[20], IN1[13], IN2);
endmodule

module UBVPPG_13_0_8 (O, IN1, IN2);
  output [21:8] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_8 U0 (O[8], IN1[0], IN2);
  UB1BPPG_1_8 U1 (O[9], IN1[1], IN2);
  UB1BPPG_2_8 U2 (O[10], IN1[2], IN2);
  UB1BPPG_3_8 U3 (O[11], IN1[3], IN2);
  UB1BPPG_4_8 U4 (O[12], IN1[4], IN2);
  UB1BPPG_5_8 U5 (O[13], IN1[5], IN2);
  UB1BPPG_6_8 U6 (O[14], IN1[6], IN2);
  UB1BPPG_7_8 U7 (O[15], IN1[7], IN2);
  UB1BPPG_8_8 U8 (O[16], IN1[8], IN2);
  UB1BPPG_9_8 U9 (O[17], IN1[9], IN2);
  UB1BPPG_10_8 U10 (O[18], IN1[10], IN2);
  UB1BPPG_11_8 U11 (O[19], IN1[11], IN2);
  UB1BPPG_12_8 U12 (O[20], IN1[12], IN2);
  UB1BPPG_13_8 U13 (O[21], IN1[13], IN2);
endmodule

module UBVPPG_13_0_9 (O, IN1, IN2);
  output [22:9] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_9 U0 (O[9], IN1[0], IN2);
  UB1BPPG_1_9 U1 (O[10], IN1[1], IN2);
  UB1BPPG_2_9 U2 (O[11], IN1[2], IN2);
  UB1BPPG_3_9 U3 (O[12], IN1[3], IN2);
  UB1BPPG_4_9 U4 (O[13], IN1[4], IN2);
  UB1BPPG_5_9 U5 (O[14], IN1[5], IN2);
  UB1BPPG_6_9 U6 (O[15], IN1[6], IN2);
  UB1BPPG_7_9 U7 (O[16], IN1[7], IN2);
  UB1BPPG_8_9 U8 (O[17], IN1[8], IN2);
  UB1BPPG_9_9 U9 (O[18], IN1[9], IN2);
  UB1BPPG_10_9 U10 (O[19], IN1[10], IN2);
  UB1BPPG_11_9 U11 (O[20], IN1[11], IN2);
  UB1BPPG_12_9 U12 (O[21], IN1[12], IN2);
  UB1BPPG_13_9 U13 (O[22], IN1[13], IN2);
endmodule

