/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: Multiplier_5_0_5_000

  Number system: Unsigned binary
  Multiplicand length: 6
  Multiplier length: 6
  Partial product generation: Simple PPG
  Partial product accumulation: Balanced delay tree
  Final stage addition: Kogge-Stone adder
----------------------------------------------------------------------------*/

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_1(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_2(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_6(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_9(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_8(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_10(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module GPGenerator(Go, Po, A, B);
  output Go;
  output Po;
  input A;
  input B;
  assign Go = A & B;
  assign Po = A ^ B;
endmodule

module CarryOperator(Go, Po, Gi1, Pi1, Gi2, Pi2);
  output Go;
  output Po;
  input Gi1;
  input Gi2;
  input Pi1;
  input Pi2;
  assign Go = Gi1 | ( Gi2 & Pi1 );
  assign Po = Pi1 & Pi2;
endmodule

module UBPriKSA_11_3(S, X, Y, Cin);
  output [12:3] S;
  input Cin;
  input [11:3] X;
  input [11:3] Y;
  wire [11:3] G0;
  wire [11:3] G1;
  wire [11:3] G2;
  wire [11:3] G3;
  wire [11:3] G4;
  wire [11:3] P0;
  wire [11:3] P1;
  wire [11:3] P2;
  wire [11:3] P3;
  wire [11:3] P4;
  assign P1[3] = P0[3];
  assign G1[3] = G0[3];
  assign P2[3] = P1[3];
  assign G2[3] = G1[3];
  assign P2[4] = P1[4];
  assign G2[4] = G1[4];
  assign P3[3] = P2[3];
  assign G3[3] = G2[3];
  assign P3[4] = P2[4];
  assign G3[4] = G2[4];
  assign P3[5] = P2[5];
  assign G3[5] = G2[5];
  assign P3[6] = P2[6];
  assign G3[6] = G2[6];
  assign P4[3] = P3[3];
  assign G4[3] = G3[3];
  assign P4[4] = P3[4];
  assign G4[4] = G3[4];
  assign P4[5] = P3[5];
  assign G4[5] = G3[5];
  assign P4[6] = P3[6];
  assign G4[6] = G3[6];
  assign P4[7] = P3[7];
  assign G4[7] = G3[7];
  assign P4[8] = P3[8];
  assign G4[8] = G3[8];
  assign P4[9] = P3[9];
  assign G4[9] = G3[9];
  assign P4[10] = P3[10];
  assign G4[10] = G3[10];
  assign S[3] = Cin ^ P0[3];
  assign S[4] = ( G4[3] | ( P4[3] & Cin ) ) ^ P0[4];
  assign S[5] = ( G4[4] | ( P4[4] & Cin ) ) ^ P0[5];
  assign S[6] = ( G4[5] | ( P4[5] & Cin ) ) ^ P0[6];
  assign S[7] = ( G4[6] | ( P4[6] & Cin ) ) ^ P0[7];
  assign S[8] = ( G4[7] | ( P4[7] & Cin ) ) ^ P0[8];
  assign S[9] = ( G4[8] | ( P4[8] & Cin ) ) ^ P0[9];
  assign S[10] = ( G4[9] | ( P4[9] & Cin ) ) ^ P0[10];
  assign S[11] = ( G4[10] | ( P4[10] & Cin ) ) ^ P0[11];
  assign S[12] = G4[11] | ( P4[11] & Cin );
  GPGenerator U0 (G0[3], P0[3], X[3], Y[3]);
  GPGenerator U1 (G0[4], P0[4], X[4], Y[4]);
  GPGenerator U2 (G0[5], P0[5], X[5], Y[5]);
  GPGenerator U3 (G0[6], P0[6], X[6], Y[6]);
  GPGenerator U4 (G0[7], P0[7], X[7], Y[7]);
  GPGenerator U5 (G0[8], P0[8], X[8], Y[8]);
  GPGenerator U6 (G0[9], P0[9], X[9], Y[9]);
  GPGenerator U7 (G0[10], P0[10], X[10], Y[10]);
  GPGenerator U8 (G0[11], P0[11], X[11], Y[11]);
  CarryOperator U9 (G1[4], P1[4], G0[4], P0[4], G0[3], P0[3]);
  CarryOperator U10 (G1[5], P1[5], G0[5], P0[5], G0[4], P0[4]);
  CarryOperator U11 (G1[6], P1[6], G0[6], P0[6], G0[5], P0[5]);
  CarryOperator U12 (G1[7], P1[7], G0[7], P0[7], G0[6], P0[6]);
  CarryOperator U13 (G1[8], P1[8], G0[8], P0[8], G0[7], P0[7]);
  CarryOperator U14 (G1[9], P1[9], G0[9], P0[9], G0[8], P0[8]);
  CarryOperator U15 (G1[10], P1[10], G0[10], P0[10], G0[9], P0[9]);
  CarryOperator U16 (G1[11], P1[11], G0[11], P0[11], G0[10], P0[10]);
  CarryOperator U17 (G2[5], P2[5], G1[5], P1[5], G1[3], P1[3]);
  CarryOperator U18 (G2[6], P2[6], G1[6], P1[6], G1[4], P1[4]);
  CarryOperator U19 (G2[7], P2[7], G1[7], P1[7], G1[5], P1[5]);
  CarryOperator U20 (G2[8], P2[8], G1[8], P1[8], G1[6], P1[6]);
  CarryOperator U21 (G2[9], P2[9], G1[9], P1[9], G1[7], P1[7]);
  CarryOperator U22 (G2[10], P2[10], G1[10], P1[10], G1[8], P1[8]);
  CarryOperator U23 (G2[11], P2[11], G1[11], P1[11], G1[9], P1[9]);
  CarryOperator U24 (G3[7], P3[7], G2[7], P2[7], G2[3], P2[3]);
  CarryOperator U25 (G3[8], P3[8], G2[8], P2[8], G2[4], P2[4]);
  CarryOperator U26 (G3[9], P3[9], G2[9], P2[9], G2[5], P2[5]);
  CarryOperator U27 (G3[10], P3[10], G2[10], P2[10], G2[6], P2[6]);
  CarryOperator U28 (G3[11], P3[11], G2[11], P2[11], G2[7], P2[7]);
  CarryOperator U29 (G4[11], P4[11], G3[11], P3[11], G3[3], P3[3]);
endmodule

module UBZero_3_3(O);
  output [3:3] O;
  assign O[3] = 0;
endmodule

module Multiplier_5_0_5_000(P, IN1, IN2);
  output [11:0] P;
  input [5:0] IN1;
  input [5:0] IN2;
  wire [12:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  MultUB_STD_BLD_KS000 U0 (W, IN1, IN2);
endmodule

module BLDCON_7_2_7_0_10000 (S1, S2, IN0, IN1, IN2, IN3);
  output [11:3] S1;
  output [11:0] S2;
  input [7:2] IN0;
  input [7:0] IN1;
  input [10:5] IN2;
  input [10:3] IN3;
  wire [11:4] W1;
  wire [10:0] W2;
  CSA_7_0_10_5_10_3 U0 (W1, W2, IN1, IN2, IN3);
  CSA_11_4_10_0_7_2 U1 (S1, S2, W1, W2, IN0);
endmodule

module BLDTR_5_0_6_1_7_2000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5);
  output [11:3] S1;
  output [11:0] S2;
  input [5:0] PP0;
  input [6:1] PP1;
  input [7:2] PP2;
  input [8:3] PP3;
  input [9:4] PP4;
  input [10:5] PP5;
  wire [7:2] W0;
  wire [7:0] W1;
  wire [10:5] W2;
  wire [10:3] W3;
  UBARYACC_5_0_6_1_000 U0 (W0, W1, PP0, PP1, PP2);
  UBARYACC_8_3_9_4_000 U1 (W2, W3, PP3, PP4, PP5);
  BLDCON_7_2_7_0_10000 U2 (S1, S2, W0, W1, W2, W3);
endmodule

module CSA_11_4_10_0_7_2 (C, S, X, Y, Z);
  output [11:3] C;
  output [11:0] S;
  input [11:4] X;
  input [10:0] Y;
  input [7:2] Z;
  UBCON_1_0 U0 (S[1:0], Y[1:0]);
  PureCSHA_3_2 U1 (C[4:3], S[3:2], Z[3:2], Y[3:2]);
  PureCSA_7_4 U2 (C[8:5], S[7:4], X[7:4], Z[7:4], Y[7:4]);
  PureCSHA_10_8 U3 (C[11:9], S[10:8], X[10:8], Y[10:8]);
  UB1DCON_11 U4 (S[11], X[11]);
endmodule

module CSA_5_0_6_1_7_2 (C, S, X, Y, Z);
  output [7:2] C;
  output [7:0] S;
  input [5:0] X;
  input [6:1] Y;
  input [7:2] Z;
  UB1DCON_0 U0 (S[0], X[0]);
  UBHA_1 U1 (C[2], S[1], Y[1], X[1]);
  PureCSA_5_2 U2 (C[6:3], S[5:2], Z[5:2], Y[5:2], X[5:2]);
  UBHA_6 U3 (C[7], S[6], Z[6], Y[6]);
  UB1DCON_7 U4 (S[7], Z[7]);
endmodule

module CSA_7_0_10_5_10_3 (C, S, X, Y, Z);
  output [11:4] C;
  output [10:0] S;
  input [7:0] X;
  input [10:5] Y;
  input [10:3] Z;
  UBCON_2_0 U0 (S[2:0], X[2:0]);
  PureCSHA_4_3 U1 (C[5:4], S[4:3], Z[4:3], X[4:3]);
  PureCSA_7_5 U2 (C[8:6], S[7:5], Y[7:5], Z[7:5], X[7:5]);
  PureCSHA_10_8 U3 (C[11:9], S[10:8], Z[10:8], Y[10:8]);
endmodule

module CSA_8_3_9_4_10_5 (C, S, X, Y, Z);
  output [10:5] C;
  output [10:3] S;
  input [8:3] X;
  input [9:4] Y;
  input [10:5] Z;
  UB1DCON_3 U0 (S[3], X[3]);
  UBHA_4 U1 (C[5], S[4], Y[4], X[4]);
  PureCSA_8_5 U2 (C[9:6], S[8:5], Z[8:5], Y[8:5], X[8:5]);
  UBHA_9 U3 (C[10], S[9], Z[9], Y[9]);
  UB1DCON_10 U4 (S[10], Z[10]);
endmodule

module MultUB_STD_BLD_KS000 (P, IN1, IN2);
  output [12:0] P;
  input [5:0] IN1;
  input [5:0] IN2;
  wire [5:0] PP0;
  wire [6:1] PP1;
  wire [7:2] PP2;
  wire [8:3] PP3;
  wire [9:4] PP4;
  wire [10:5] PP5;
  wire [11:3] S1;
  wire [11:0] S2;
  UBPPG_5_0_5_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, IN1, IN2);
  BLDTR_5_0_6_1_7_2000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5);
  UBKSA_11_3_11_0 U2 (P, S1, S2);
endmodule

module PureCSA_5_2 (C, S, X, Y, Z);
  output [6:3] C;
  output [5:2] S;
  input [5:2] X;
  input [5:2] Y;
  input [5:2] Z;
  UBFA_2 U0 (C[3], S[2], X[2], Y[2], Z[2]);
  UBFA_3 U1 (C[4], S[3], X[3], Y[3], Z[3]);
  UBFA_4 U2 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U3 (C[6], S[5], X[5], Y[5], Z[5]);
endmodule

module PureCSA_7_4 (C, S, X, Y, Z);
  output [8:5] C;
  output [7:4] S;
  input [7:4] X;
  input [7:4] Y;
  input [7:4] Z;
  UBFA_4 U0 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U1 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U2 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U3 (C[8], S[7], X[7], Y[7], Z[7]);
endmodule

module PureCSA_7_5 (C, S, X, Y, Z);
  output [8:6] C;
  output [7:5] S;
  input [7:5] X;
  input [7:5] Y;
  input [7:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
endmodule

module PureCSA_8_5 (C, S, X, Y, Z);
  output [9:6] C;
  output [8:5] S;
  input [8:5] X;
  input [8:5] Y;
  input [8:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U3 (C[9], S[8], X[8], Y[8], Z[8]);
endmodule

module PureCSHA_10_8 (C, S, X, Y);
  output [11:9] C;
  output [10:8] S;
  input [10:8] X;
  input [10:8] Y;
  UBHA_8 U0 (C[9], S[8], X[8], Y[8]);
  UBHA_9 U1 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U2 (C[11], S[10], X[10], Y[10]);
endmodule

module PureCSHA_3_2 (C, S, X, Y);
  output [4:3] C;
  output [3:2] S;
  input [3:2] X;
  input [3:2] Y;
  UBHA_2 U0 (C[3], S[2], X[2], Y[2]);
  UBHA_3 U1 (C[4], S[3], X[3], Y[3]);
endmodule

module PureCSHA_4_3 (C, S, X, Y);
  output [5:4] C;
  output [4:3] S;
  input [4:3] X;
  input [4:3] Y;
  UBHA_3 U0 (C[4], S[3], X[3], Y[3]);
  UBHA_4 U1 (C[5], S[4], X[4], Y[4]);
endmodule

module UBARYACC_5_0_6_1_000 (S1, S2, PP0, PP1, PP2);
  output [7:2] S1;
  output [7:0] S2;
  input [5:0] PP0;
  input [6:1] PP1;
  input [7:2] PP2;
  CSA_5_0_6_1_7_2 U0 (S1, S2, PP0, PP1, PP2);
endmodule

module UBARYACC_8_3_9_4_000 (S1, S2, PP0, PP1, PP2);
  output [10:5] S1;
  output [10:3] S2;
  input [8:3] PP0;
  input [9:4] PP1;
  input [10:5] PP2;
  CSA_8_3_9_4_10_5 U0 (S1, S2, PP0, PP1, PP2);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBKSA_11_3_11_0 (S, X, Y);
  output [12:0] S;
  input [11:3] X;
  input [11:0] Y;
  UBPureKSA_11_3 U0 (S[12:3], X[11:3], Y[11:3]);
  UBCON_2_0 U1 (S[2:0], Y[2:0]);
endmodule

module UBPPG_5_0_5_0 (PP0, PP1, PP2, PP3, PP4, PP5, IN1, IN2);
  output [5:0] PP0;
  output [6:1] PP1;
  output [7:2] PP2;
  output [8:3] PP3;
  output [9:4] PP4;
  output [10:5] PP5;
  input [5:0] IN1;
  input [5:0] IN2;
  UBVPPG_5_0_0 U0 (PP0, IN1, IN2[0]);
  UBVPPG_5_0_1 U1 (PP1, IN1, IN2[1]);
  UBVPPG_5_0_2 U2 (PP2, IN1, IN2[2]);
  UBVPPG_5_0_3 U3 (PP3, IN1, IN2[3]);
  UBVPPG_5_0_4 U4 (PP4, IN1, IN2[4]);
  UBVPPG_5_0_5 U5 (PP5, IN1, IN2[5]);
endmodule

module UBPureKSA_11_3 (S, X, Y);
  output [12:3] S;
  input [11:3] X;
  input [11:3] Y;
  wire C;
  UBPriKSA_11_3 U0 (S, X, Y, C);
  UBZero_3_3 U1 (C);
endmodule

module UBVPPG_5_0_0 (O, IN1, IN2);
  output [5:0] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
endmodule

module UBVPPG_5_0_1 (O, IN1, IN2);
  output [6:1] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_1 U0 (O[1], IN1[0], IN2);
  UB1BPPG_1_1 U1 (O[2], IN1[1], IN2);
  UB1BPPG_2_1 U2 (O[3], IN1[2], IN2);
  UB1BPPG_3_1 U3 (O[4], IN1[3], IN2);
  UB1BPPG_4_1 U4 (O[5], IN1[4], IN2);
  UB1BPPG_5_1 U5 (O[6], IN1[5], IN2);
endmodule

module UBVPPG_5_0_2 (O, IN1, IN2);
  output [7:2] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
endmodule

module UBVPPG_5_0_3 (O, IN1, IN2);
  output [8:3] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_3 U0 (O[3], IN1[0], IN2);
  UB1BPPG_1_3 U1 (O[4], IN1[1], IN2);
  UB1BPPG_2_3 U2 (O[5], IN1[2], IN2);
  UB1BPPG_3_3 U3 (O[6], IN1[3], IN2);
  UB1BPPG_4_3 U4 (O[7], IN1[4], IN2);
  UB1BPPG_5_3 U5 (O[8], IN1[5], IN2);
endmodule

module UBVPPG_5_0_4 (O, IN1, IN2);
  output [9:4] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
endmodule

module UBVPPG_5_0_5 (O, IN1, IN2);
  output [10:5] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_5 U0 (O[5], IN1[0], IN2);
  UB1BPPG_1_5 U1 (O[6], IN1[1], IN2);
  UB1BPPG_2_5 U2 (O[7], IN1[2], IN2);
  UB1BPPG_3_5 U3 (O[8], IN1[3], IN2);
  UB1BPPG_4_5 U4 (O[9], IN1[4], IN2);
  UB1BPPG_5_5 U5 (O[10], IN1[5], IN2);
endmodule

