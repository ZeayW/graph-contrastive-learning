/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: Multiplier_9_0_9_000

  Number system: Unsigned binary
  Multiplicand length: 10
  Multiplier length: 10
  Partial product generation: Simple PPG
  Partial product accumulation: Dadda tree
  Final stage addition: Ripple carry adder
----------------------------------------------------------------------------*/

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UBHA_9(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_10(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_6(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_7(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_8(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_12(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_13(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_5(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_14(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_15(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_16(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_17(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_1(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_2(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_18(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBZero_1_1(O);
  output [1:1] O;
  assign O[1] = 0;
endmodule

module Multiplier_9_0_9_000(P, IN1, IN2);
  output [19:0] P;
  input [9:0] IN1;
  input [9:0] IN2;
  wire [19:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  assign P[12] = W[12];
  assign P[13] = W[13];
  assign P[14] = W[14];
  assign P[15] = W[15];
  assign P[16] = W[16];
  assign P[17] = W[17];
  assign P[18] = W[18];
  assign P[19] = W[19];
  MultUB_STD_DAD_RC000 U0 (W, IN1, IN2);
endmodule

module DADTR_18_0_17_1_1000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8);
  output [18:0] S1;
  output [18:1] S2;
  input [18:0] PP0;
  input [17:1] PP1;
  input [16:2] PP2;
  input [15:3] PP3;
  input [14:4] PP4;
  input [13:5] PP5;
  input [12:6] PP6;
  input [11:7] PP7;
  input [11:8] PP8;
  wire [18:0] W0;
  wire [17:1] W1;
  wire [16:2] W2;
  wire [15:3] W3;
  wire [14:4] W4;
  wire [14:5] W5;
  UBHA_6 U0 (W3[7], W5[6], PP0[6], PP1[6]);
  UBFA_7 U1 (W1[8], W4[7], PP0[7], PP1[7], PP2[7]);
  UBHA_7 U2 (W2[8], W5[7], PP3[7], PP4[7]);
  UBFA_8 U3 (W0[9], W3[8], PP0[8], PP1[8], PP2[8]);
  UBFA_8 U4 (W1[9], W4[8], PP3[8], PP4[8], PP5[8]);
  UBHA_8 U5 (W2[9], W5[8], PP6[8], PP7[8]);
  UBFA_9 U6 (W0[10], W3[9], PP0[9], PP1[9], PP2[9]);
  UBFA_9 U7 (W1[10], W4[9], PP3[9], PP4[9], PP5[9]);
  UBFA_9 U8 (W2[10], W5[9], PP6[9], PP7[9], PP8[9]);
  UBFA_10 U9 (W0[11], W3[10], PP0[10], PP1[10], PP2[10]);
  UBFA_10 U10 (W1[11], W4[10], PP3[10], PP4[10], PP5[10]);
  UBFA_10 U11 (W2[11], W5[10], PP6[10], PP7[10], PP8[10]);
  UBFA_11 U12 (W1[12], W3[11], PP0[11], PP1[11], PP2[11]);
  UBFA_11 U13 (W2[12], W4[11], PP3[11], PP4[11], PP5[11]);
  UBFA_11 U14 (W3[12], W5[11], PP6[11], PP7[11], PP8[11]);
  UBFA_12 U15 (W3[13], W4[12], PP0[12], PP1[12], PP2[12]);
  UBFA_12 U16 (W4[13], W5[12], PP3[12], PP4[12], PP5[12]);
  UBFA_13 U17 (W5[14], W5[13], PP0[13], PP1[13], PP2[13]);
  UBCON_5_0 U18 (W0[5:0], PP0[5:0]);
  UB1DCON_6 U19 (W0[6], PP2[6]);
  UB1DCON_7 U20 (W0[7], PP5[7]);
  UB1DCON_8 U21 (W0[8], PP8[8]);
  UB1DCON_12 U22 (W0[12], PP6[12]);
  UB1DCON_13 U23 (W0[13], PP3[13]);
  UBCON_18_14 U24 (W0[18:14], PP0[18:14]);
  UBCON_5_1 U25 (W1[5:1], PP1[5:1]);
  UB1DCON_6 U26 (W1[6], PP3[6]);
  UB1DCON_7 U27 (W1[7], PP6[7]);
  UB1DCON_13 U28 (W1[13], PP4[13]);
  UBCON_17_14 U29 (W1[17:14], PP1[17:14]);
  UBCON_5_2 U30 (W2[5:2], PP2[5:2]);
  UB1DCON_6 U31 (W2[6], PP4[6]);
  UB1DCON_7 U32 (W2[7], PP7[7]);
  UB1DCON_13 U33 (W2[13], PP5[13]);
  UBCON_16_14 U34 (W2[16:14], PP2[16:14]);
  UBCON_5_3 U35 (W3[5:3], PP3[5:3]);
  UB1DCON_6 U36 (W3[6], PP5[6]);
  UBCON_15_14 U37 (W3[15:14], PP3[15:14]);
  UBCON_5_4 U38 (W4[5:4], PP4[5:4]);
  UB1DCON_6 U39 (W4[6], PP6[6]);
  UB1DCON_14 U40 (W4[14], PP4[14]);
  UB1DCON_5 U41 (W5[5], PP5[5]);
  DADTR_18_0_17_1_1001 U42 (S1, S2, W0, W1, W2, W3, W4, W5);
endmodule

module DADTR_18_0_17_1_1001 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5);
  output [18:0] S1;
  output [18:1] S2;
  input [18:0] PP0;
  input [17:1] PP1;
  input [16:2] PP2;
  input [15:3] PP3;
  input [14:4] PP4;
  input [14:5] PP5;
  wire [18:0] W0;
  wire [17:1] W1;
  wire [16:2] W2;
  wire [16:3] W3;
  UBHA_4 U0 (W1[5], W3[4], PP0[4], PP1[4]);
  UBFA_5 U1 (W0[6], W2[5], PP0[5], PP1[5], PP2[5]);
  UBHA_5 U2 (W1[6], W3[5], PP3[5], PP4[5]);
  UBFA_6 U3 (W0[7], W2[6], PP0[6], PP1[6], PP2[6]);
  UBFA_6 U4 (W1[7], W3[6], PP3[6], PP4[6], PP5[6]);
  UBFA_7 U5 (W0[8], W2[7], PP0[7], PP1[7], PP2[7]);
  UBFA_7 U6 (W1[8], W3[7], PP3[7], PP4[7], PP5[7]);
  UBFA_8 U7 (W0[9], W2[8], PP0[8], PP1[8], PP2[8]);
  UBFA_8 U8 (W1[9], W3[8], PP3[8], PP4[8], PP5[8]);
  UBFA_9 U9 (W0[10], W2[9], PP0[9], PP1[9], PP2[9]);
  UBFA_9 U10 (W1[10], W3[9], PP3[9], PP4[9], PP5[9]);
  UBFA_10 U11 (W0[11], W2[10], PP0[10], PP1[10], PP2[10]);
  UBFA_10 U12 (W1[11], W3[10], PP3[10], PP4[10], PP5[10]);
  UBFA_11 U13 (W0[12], W2[11], PP0[11], PP1[11], PP2[11]);
  UBFA_11 U14 (W1[12], W3[11], PP3[11], PP4[11], PP5[11]);
  UBFA_12 U15 (W0[13], W2[12], PP0[12], PP1[12], PP2[12]);
  UBFA_12 U16 (W1[13], W3[12], PP3[12], PP4[12], PP5[12]);
  UBFA_13 U17 (W0[14], W2[13], PP0[13], PP1[13], PP2[13]);
  UBFA_13 U18 (W1[14], W3[13], PP3[13], PP4[13], PP5[13]);
  UBFA_14 U19 (W1[15], W2[14], PP0[14], PP1[14], PP2[14]);
  UBFA_14 U20 (W2[15], W3[14], PP3[14], PP4[14], PP5[14]);
  UBFA_15 U21 (W3[16], W3[15], PP0[15], PP1[15], PP2[15]);
  UBCON_3_0 U22 (W0[3:0], PP0[3:0]);
  UB1DCON_4 U23 (W0[4], PP2[4]);
  UB1DCON_5 U24 (W0[5], PP5[5]);
  UB1DCON_15 U25 (W0[15], PP3[15]);
  UBCON_18_16 U26 (W0[18:16], PP0[18:16]);
  UBCON_3_1 U27 (W1[3:1], PP1[3:1]);
  UB1DCON_4 U28 (W1[4], PP3[4]);
  UBCON_17_16 U29 (W1[17:16], PP1[17:16]);
  UBCON_3_2 U30 (W2[3:2], PP2[3:2]);
  UB1DCON_4 U31 (W2[4], PP4[4]);
  UB1DCON_16 U32 (W2[16], PP2[16]);
  UB1DCON_3 U33 (W3[3], PP3[3]);
  DADTR_18_0_17_1_1002 U34 (S1, S2, W0, W1, W2, W3);
endmodule

module DADTR_18_0_17_1_1002 (S1, S2, PP0, PP1, PP2, PP3);
  output [18:0] S1;
  output [18:1] S2;
  input [18:0] PP0;
  input [17:1] PP1;
  input [16:2] PP2;
  input [16:3] PP3;
  wire [18:0] W0;
  wire [17:1] W1;
  wire [17:2] W2;
  UBHA_3 U0 (W1[4], W2[3], PP0[3], PP1[3]);
  UBFA_4 U1 (W1[5], W2[4], PP0[4], PP1[4], PP2[4]);
  UBFA_5 U2 (W1[6], W2[5], PP0[5], PP1[5], PP2[5]);
  UBFA_6 U3 (W1[7], W2[6], PP0[6], PP1[6], PP2[6]);
  UBFA_7 U4 (W1[8], W2[7], PP0[7], PP1[7], PP2[7]);
  UBFA_8 U5 (W1[9], W2[8], PP0[8], PP1[8], PP2[8]);
  UBFA_9 U6 (W1[10], W2[9], PP0[9], PP1[9], PP2[9]);
  UBFA_10 U7 (W1[11], W2[10], PP0[10], PP1[10], PP2[10]);
  UBFA_11 U8 (W1[12], W2[11], PP0[11], PP1[11], PP2[11]);
  UBFA_12 U9 (W1[13], W2[12], PP0[12], PP1[12], PP2[12]);
  UBFA_13 U10 (W1[14], W2[13], PP0[13], PP1[13], PP2[13]);
  UBFA_14 U11 (W1[15], W2[14], PP0[14], PP1[14], PP2[14]);
  UBFA_15 U12 (W1[16], W2[15], PP0[15], PP1[15], PP2[15]);
  UBFA_16 U13 (W2[17], W2[16], PP0[16], PP1[16], PP2[16]);
  UBCON_2_0 U14 (W0[2:0], PP0[2:0]);
  UB1DCON_3 U15 (W0[3], PP2[3]);
  UBCON_16_4 U16 (W0[16:4], PP3[16:4]);
  UBCON_18_17 U17 (W0[18:17], PP0[18:17]);
  UBCON_2_1 U18 (W1[2:1], PP1[2:1]);
  UB1DCON_3 U19 (W1[3], PP3[3]);
  UB1DCON_17 U20 (W1[17], PP1[17]);
  UB1DCON_2 U21 (W2[2], PP2[2]);
  DADTR_18_0_17_1_1003 U22 (S1, S2, W0, W1, W2);
endmodule

module DADTR_18_0_17_1_1003 (S1, S2, PP0, PP1, PP2);
  output [18:0] S1;
  output [18:1] S2;
  input [18:0] PP0;
  input [17:1] PP1;
  input [17:2] PP2;
  wire [18:0] W0;
  wire [18:1] W1;
  UBHA_2 U0 (W0[3], W1[2], PP0[2], PP1[2]);
  UBFA_3 U1 (W0[4], W1[3], PP0[3], PP1[3], PP2[3]);
  UBFA_4 U2 (W0[5], W1[4], PP0[4], PP1[4], PP2[4]);
  UBFA_5 U3 (W0[6], W1[5], PP0[5], PP1[5], PP2[5]);
  UBFA_6 U4 (W0[7], W1[6], PP0[6], PP1[6], PP2[6]);
  UBFA_7 U5 (W0[8], W1[7], PP0[7], PP1[7], PP2[7]);
  UBFA_8 U6 (W0[9], W1[8], PP0[8], PP1[8], PP2[8]);
  UBFA_9 U7 (W0[10], W1[9], PP0[9], PP1[9], PP2[9]);
  UBFA_10 U8 (W0[11], W1[10], PP0[10], PP1[10], PP2[10]);
  UBFA_11 U9 (W0[12], W1[11], PP0[11], PP1[11], PP2[11]);
  UBFA_12 U10 (W0[13], W1[12], PP0[12], PP1[12], PP2[12]);
  UBFA_13 U11 (W0[14], W1[13], PP0[13], PP1[13], PP2[13]);
  UBFA_14 U12 (W0[15], W1[14], PP0[14], PP1[14], PP2[14]);
  UBFA_15 U13 (W0[16], W1[15], PP0[15], PP1[15], PP2[15]);
  UBFA_16 U14 (W0[17], W1[16], PP0[16], PP1[16], PP2[16]);
  UBFA_17 U15 (W1[18], W1[17], PP0[17], PP1[17], PP2[17]);
  UBCON_1_0 U16 (W0[1:0], PP0[1:0]);
  UB1DCON_2 U17 (W0[2], PP2[2]);
  UB1DCON_18 U18 (W0[18], PP0[18]);
  UB1DCON_1 U19 (W1[1], PP1[1]);
  DADTR_18_0_18_1 U20 (S1, S2, W0, W1);
endmodule

module DADTR_18_0_18_1 (S1, S2, PP0, PP1);
  output [18:0] S1;
  output [18:1] S2;
  input [18:0] PP0;
  input [18:1] PP1;
  UBCON_18_0 U0 (S1, PP0);
  UBCON_18_1 U1 (S2, PP1);
endmodule

module DADTR_9_0_10_1_11000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9);
  output [18:0] S1;
  output [18:1] S2;
  input [9:0] PP0;
  input [10:1] PP1;
  input [11:2] PP2;
  input [12:3] PP3;
  input [13:4] PP4;
  input [14:5] PP5;
  input [15:6] PP6;
  input [16:7] PP7;
  input [17:8] PP8;
  input [18:9] PP9;
  wire [18:0] W0;
  wire [17:1] W1;
  wire [16:2] W2;
  wire [15:3] W3;
  wire [14:4] W4;
  wire [13:5] W5;
  wire [12:6] W6;
  wire [11:7] W7;
  wire [11:8] W8;
  UBHA_9 U0 (W7[10], W8[9], PP0[9], PP1[9]);
  UBHA_10 U1 (W8[11], W8[10], PP1[10], PP2[10]);
  UBCON_8_0 U2 (W0[8:0], PP0[8:0]);
  UB1DCON_9 U3 (W0[9], PP2[9]);
  UB1DCON_10 U4 (W0[10], PP3[10]);
  UB1DCON_11 U5 (W0[11], PP2[11]);
  UB1DCON_12 U6 (W0[12], PP3[12]);
  UB1DCON_13 U7 (W0[13], PP4[13]);
  UB1DCON_14 U8 (W0[14], PP5[14]);
  UB1DCON_15 U9 (W0[15], PP6[15]);
  UB1DCON_16 U10 (W0[16], PP7[16]);
  UB1DCON_17 U11 (W0[17], PP8[17]);
  UB1DCON_18 U12 (W0[18], PP9[18]);
  UBCON_8_1 U13 (W1[8:1], PP1[8:1]);
  UB1DCON_9 U14 (W1[9], PP3[9]);
  UB1DCON_10 U15 (W1[10], PP4[10]);
  UB1DCON_11 U16 (W1[11], PP3[11]);
  UB1DCON_12 U17 (W1[12], PP4[12]);
  UB1DCON_13 U18 (W1[13], PP5[13]);
  UB1DCON_14 U19 (W1[14], PP6[14]);
  UB1DCON_15 U20 (W1[15], PP7[15]);
  UB1DCON_16 U21 (W1[16], PP8[16]);
  UB1DCON_17 U22 (W1[17], PP9[17]);
  UBCON_8_2 U23 (W2[8:2], PP2[8:2]);
  UB1DCON_9 U24 (W2[9], PP4[9]);
  UB1DCON_10 U25 (W2[10], PP5[10]);
  UB1DCON_11 U26 (W2[11], PP4[11]);
  UB1DCON_12 U27 (W2[12], PP5[12]);
  UB1DCON_13 U28 (W2[13], PP6[13]);
  UB1DCON_14 U29 (W2[14], PP7[14]);
  UB1DCON_15 U30 (W2[15], PP8[15]);
  UB1DCON_16 U31 (W2[16], PP9[16]);
  UBCON_8_3 U32 (W3[8:3], PP3[8:3]);
  UB1DCON_9 U33 (W3[9], PP5[9]);
  UB1DCON_10 U34 (W3[10], PP6[10]);
  UB1DCON_11 U35 (W3[11], PP5[11]);
  UB1DCON_12 U36 (W3[12], PP6[12]);
  UB1DCON_13 U37 (W3[13], PP7[13]);
  UB1DCON_14 U38 (W3[14], PP8[14]);
  UB1DCON_15 U39 (W3[15], PP9[15]);
  UBCON_8_4 U40 (W4[8:4], PP4[8:4]);
  UB1DCON_9 U41 (W4[9], PP6[9]);
  UB1DCON_10 U42 (W4[10], PP7[10]);
  UB1DCON_11 U43 (W4[11], PP6[11]);
  UB1DCON_12 U44 (W4[12], PP7[12]);
  UB1DCON_13 U45 (W4[13], PP8[13]);
  UB1DCON_14 U46 (W4[14], PP9[14]);
  UBCON_8_5 U47 (W5[8:5], PP5[8:5]);
  UB1DCON_9 U48 (W5[9], PP7[9]);
  UB1DCON_10 U49 (W5[10], PP8[10]);
  UB1DCON_11 U50 (W5[11], PP7[11]);
  UB1DCON_12 U51 (W5[12], PP8[12]);
  UB1DCON_13 U52 (W5[13], PP9[13]);
  UBCON_8_6 U53 (W6[8:6], PP6[8:6]);
  UB1DCON_9 U54 (W6[9], PP8[9]);
  UB1DCON_10 U55 (W6[10], PP9[10]);
  UB1DCON_11 U56 (W6[11], PP8[11]);
  UB1DCON_12 U57 (W6[12], PP9[12]);
  UBCON_8_7 U58 (W7[8:7], PP7[8:7]);
  UB1DCON_9 U59 (W7[9], PP9[9]);
  UB1DCON_11 U60 (W7[11], PP9[11]);
  UB1DCON_8 U61 (W8[8], PP8[8]);
  DADTR_18_0_17_1_1000 U62 (S1, S2, W0, W1, W2, W3, W4, W5, W6, W7, W8);
endmodule

module MultUB_STD_DAD_RC000 (P, IN1, IN2);
  output [19:0] P;
  input [9:0] IN1;
  input [9:0] IN2;
  wire [9:0] PP0;
  wire [10:1] PP1;
  wire [11:2] PP2;
  wire [12:3] PP3;
  wire [13:4] PP4;
  wire [14:5] PP5;
  wire [15:6] PP6;
  wire [16:7] PP7;
  wire [17:8] PP8;
  wire [18:9] PP9;
  wire [18:0] S1;
  wire [18:1] S2;
  UBPPG_9_0_9_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, IN1, IN2);
  DADTR_9_0_10_1_11000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9);
  UBRCA_18_0_18_1 U2 (P, S1, S2);
endmodule

module UBCON_15_14 (O, I);
  output [15:14] O;
  input [15:14] I;
  UB1DCON_14 U0 (O[14], I[14]);
  UB1DCON_15 U1 (O[15], I[15]);
endmodule

module UBCON_16_14 (O, I);
  output [16:14] O;
  input [16:14] I;
  UB1DCON_14 U0 (O[14], I[14]);
  UB1DCON_15 U1 (O[15], I[15]);
  UB1DCON_16 U2 (O[16], I[16]);
endmodule

module UBCON_16_4 (O, I);
  output [16:4] O;
  input [16:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
  UB1DCON_11 U7 (O[11], I[11]);
  UB1DCON_12 U8 (O[12], I[12]);
  UB1DCON_13 U9 (O[13], I[13]);
  UB1DCON_14 U10 (O[14], I[14]);
  UB1DCON_15 U11 (O[15], I[15]);
  UB1DCON_16 U12 (O[16], I[16]);
endmodule

module UBCON_17_14 (O, I);
  output [17:14] O;
  input [17:14] I;
  UB1DCON_14 U0 (O[14], I[14]);
  UB1DCON_15 U1 (O[15], I[15]);
  UB1DCON_16 U2 (O[16], I[16]);
  UB1DCON_17 U3 (O[17], I[17]);
endmodule

module UBCON_17_16 (O, I);
  output [17:16] O;
  input [17:16] I;
  UB1DCON_16 U0 (O[16], I[16]);
  UB1DCON_17 U1 (O[17], I[17]);
endmodule

module UBCON_18_0 (O, I);
  output [18:0] O;
  input [18:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
  UB1DCON_13 U13 (O[13], I[13]);
  UB1DCON_14 U14 (O[14], I[14]);
  UB1DCON_15 U15 (O[15], I[15]);
  UB1DCON_16 U16 (O[16], I[16]);
  UB1DCON_17 U17 (O[17], I[17]);
  UB1DCON_18 U18 (O[18], I[18]);
endmodule

module UBCON_18_1 (O, I);
  output [18:1] O;
  input [18:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
  UB1DCON_6 U5 (O[6], I[6]);
  UB1DCON_7 U6 (O[7], I[7]);
  UB1DCON_8 U7 (O[8], I[8]);
  UB1DCON_9 U8 (O[9], I[9]);
  UB1DCON_10 U9 (O[10], I[10]);
  UB1DCON_11 U10 (O[11], I[11]);
  UB1DCON_12 U11 (O[12], I[12]);
  UB1DCON_13 U12 (O[13], I[13]);
  UB1DCON_14 U13 (O[14], I[14]);
  UB1DCON_15 U14 (O[15], I[15]);
  UB1DCON_16 U15 (O[16], I[16]);
  UB1DCON_17 U16 (O[17], I[17]);
  UB1DCON_18 U17 (O[18], I[18]);
endmodule

module UBCON_18_14 (O, I);
  output [18:14] O;
  input [18:14] I;
  UB1DCON_14 U0 (O[14], I[14]);
  UB1DCON_15 U1 (O[15], I[15]);
  UB1DCON_16 U2 (O[16], I[16]);
  UB1DCON_17 U3 (O[17], I[17]);
  UB1DCON_18 U4 (O[18], I[18]);
endmodule

module UBCON_18_16 (O, I);
  output [18:16] O;
  input [18:16] I;
  UB1DCON_16 U0 (O[16], I[16]);
  UB1DCON_17 U1 (O[17], I[17]);
  UB1DCON_18 U2 (O[18], I[18]);
endmodule

module UBCON_18_17 (O, I);
  output [18:17] O;
  input [18:17] I;
  UB1DCON_17 U0 (O[17], I[17]);
  UB1DCON_18 U1 (O[18], I[18]);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBCON_2_1 (O, I);
  output [2:1] O;
  input [2:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
endmodule

module UBCON_3_0 (O, I);
  output [3:0] O;
  input [3:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
endmodule

module UBCON_3_1 (O, I);
  output [3:1] O;
  input [3:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
endmodule

module UBCON_3_2 (O, I);
  output [3:2] O;
  input [3:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
endmodule

module UBCON_5_0 (O, I);
  output [5:0] O;
  input [5:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
endmodule

module UBCON_5_1 (O, I);
  output [5:1] O;
  input [5:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
endmodule

module UBCON_5_2 (O, I);
  output [5:2] O;
  input [5:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
endmodule

module UBCON_5_3 (O, I);
  output [5:3] O;
  input [5:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
endmodule

module UBCON_5_4 (O, I);
  output [5:4] O;
  input [5:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
endmodule

module UBCON_8_0 (O, I);
  output [8:0] O;
  input [8:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
endmodule

module UBCON_8_1 (O, I);
  output [8:1] O;
  input [8:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
  UB1DCON_6 U5 (O[6], I[6]);
  UB1DCON_7 U6 (O[7], I[7]);
  UB1DCON_8 U7 (O[8], I[8]);
endmodule

module UBCON_8_2 (O, I);
  output [8:2] O;
  input [8:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
  UB1DCON_6 U4 (O[6], I[6]);
  UB1DCON_7 U5 (O[7], I[7]);
  UB1DCON_8 U6 (O[8], I[8]);
endmodule

module UBCON_8_3 (O, I);
  output [8:3] O;
  input [8:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
  UB1DCON_6 U3 (O[6], I[6]);
  UB1DCON_7 U4 (O[7], I[7]);
  UB1DCON_8 U5 (O[8], I[8]);
endmodule

module UBCON_8_4 (O, I);
  output [8:4] O;
  input [8:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
endmodule

module UBCON_8_5 (O, I);
  output [8:5] O;
  input [8:5] I;
  UB1DCON_5 U0 (O[5], I[5]);
  UB1DCON_6 U1 (O[6], I[6]);
  UB1DCON_7 U2 (O[7], I[7]);
  UB1DCON_8 U3 (O[8], I[8]);
endmodule

module UBCON_8_6 (O, I);
  output [8:6] O;
  input [8:6] I;
  UB1DCON_6 U0 (O[6], I[6]);
  UB1DCON_7 U1 (O[7], I[7]);
  UB1DCON_8 U2 (O[8], I[8]);
endmodule

module UBCON_8_7 (O, I);
  output [8:7] O;
  input [8:7] I;
  UB1DCON_7 U0 (O[7], I[7]);
  UB1DCON_8 U1 (O[8], I[8]);
endmodule

module UBPPG_9_0_9_0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, IN1, IN2);
  output [9:0] PP0;
  output [10:1] PP1;
  output [11:2] PP2;
  output [12:3] PP3;
  output [13:4] PP4;
  output [14:5] PP5;
  output [15:6] PP6;
  output [16:7] PP7;
  output [17:8] PP8;
  output [18:9] PP9;
  input [9:0] IN1;
  input [9:0] IN2;
  UBVPPG_9_0_0 U0 (PP0, IN1, IN2[0]);
  UBVPPG_9_0_1 U1 (PP1, IN1, IN2[1]);
  UBVPPG_9_0_2 U2 (PP2, IN1, IN2[2]);
  UBVPPG_9_0_3 U3 (PP3, IN1, IN2[3]);
  UBVPPG_9_0_4 U4 (PP4, IN1, IN2[4]);
  UBVPPG_9_0_5 U5 (PP5, IN1, IN2[5]);
  UBVPPG_9_0_6 U6 (PP6, IN1, IN2[6]);
  UBVPPG_9_0_7 U7 (PP7, IN1, IN2[7]);
  UBVPPG_9_0_8 U8 (PP8, IN1, IN2[8]);
  UBVPPG_9_0_9 U9 (PP9, IN1, IN2[9]);
endmodule

module UBPriRCA_18_1 (S, X, Y, Cin);
  output [19:1] S;
  input Cin;
  input [18:1] X;
  input [18:1] Y;
  wire C10;
  wire C11;
  wire C12;
  wire C13;
  wire C14;
  wire C15;
  wire C16;
  wire C17;
  wire C18;
  wire C2;
  wire C3;
  wire C4;
  wire C5;
  wire C6;
  wire C7;
  wire C8;
  wire C9;
  UBFA_1 U0 (C2, S[1], X[1], Y[1], Cin);
  UBFA_2 U1 (C3, S[2], X[2], Y[2], C2);
  UBFA_3 U2 (C4, S[3], X[3], Y[3], C3);
  UBFA_4 U3 (C5, S[4], X[4], Y[4], C4);
  UBFA_5 U4 (C6, S[5], X[5], Y[5], C5);
  UBFA_6 U5 (C7, S[6], X[6], Y[6], C6);
  UBFA_7 U6 (C8, S[7], X[7], Y[7], C7);
  UBFA_8 U7 (C9, S[8], X[8], Y[8], C8);
  UBFA_9 U8 (C10, S[9], X[9], Y[9], C9);
  UBFA_10 U9 (C11, S[10], X[10], Y[10], C10);
  UBFA_11 U10 (C12, S[11], X[11], Y[11], C11);
  UBFA_12 U11 (C13, S[12], X[12], Y[12], C12);
  UBFA_13 U12 (C14, S[13], X[13], Y[13], C13);
  UBFA_14 U13 (C15, S[14], X[14], Y[14], C14);
  UBFA_15 U14 (C16, S[15], X[15], Y[15], C15);
  UBFA_16 U15 (C17, S[16], X[16], Y[16], C16);
  UBFA_17 U16 (C18, S[17], X[17], Y[17], C17);
  UBFA_18 U17 (S[19], S[18], X[18], Y[18], C18);
endmodule

module UBPureRCA_18_1 (S, X, Y);
  output [19:1] S;
  input [18:1] X;
  input [18:1] Y;
  wire C;
  UBPriRCA_18_1 U0 (S, X, Y, C);
  UBZero_1_1 U1 (C);
endmodule

module UBRCA_18_0_18_1 (S, X, Y);
  output [19:0] S;
  input [18:0] X;
  input [18:1] Y;
  UBPureRCA_18_1 U0 (S[19:1], X[18:1], Y[18:1]);
  UB1DCON_0 U1 (S[0], X[0]);
endmodule

module UBVPPG_9_0_0 (O, IN1, IN2);
  output [9:0] O;
  input [9:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
  UB1BPPG_6_0 U6 (O[6], IN1[6], IN2);
  UB1BPPG_7_0 U7 (O[7], IN1[7], IN2);
  UB1BPPG_8_0 U8 (O[8], IN1[8], IN2);
  UB1BPPG_9_0 U9 (O[9], IN1[9], IN2);
endmodule

module UBVPPG_9_0_1 (O, IN1, IN2);
  output [10:1] O;
  input [9:0] IN1;
  input IN2;
  UB1BPPG_0_1 U0 (O[1], IN1[0], IN2);
  UB1BPPG_1_1 U1 (O[2], IN1[1], IN2);
  UB1BPPG_2_1 U2 (O[3], IN1[2], IN2);
  UB1BPPG_3_1 U3 (O[4], IN1[3], IN2);
  UB1BPPG_4_1 U4 (O[5], IN1[4], IN2);
  UB1BPPG_5_1 U5 (O[6], IN1[5], IN2);
  UB1BPPG_6_1 U6 (O[7], IN1[6], IN2);
  UB1BPPG_7_1 U7 (O[8], IN1[7], IN2);
  UB1BPPG_8_1 U8 (O[9], IN1[8], IN2);
  UB1BPPG_9_1 U9 (O[10], IN1[9], IN2);
endmodule

module UBVPPG_9_0_2 (O, IN1, IN2);
  output [11:2] O;
  input [9:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
  UB1BPPG_6_2 U6 (O[8], IN1[6], IN2);
  UB1BPPG_7_2 U7 (O[9], IN1[7], IN2);
  UB1BPPG_8_2 U8 (O[10], IN1[8], IN2);
  UB1BPPG_9_2 U9 (O[11], IN1[9], IN2);
endmodule

module UBVPPG_9_0_3 (O, IN1, IN2);
  output [12:3] O;
  input [9:0] IN1;
  input IN2;
  UB1BPPG_0_3 U0 (O[3], IN1[0], IN2);
  UB1BPPG_1_3 U1 (O[4], IN1[1], IN2);
  UB1BPPG_2_3 U2 (O[5], IN1[2], IN2);
  UB1BPPG_3_3 U3 (O[6], IN1[3], IN2);
  UB1BPPG_4_3 U4 (O[7], IN1[4], IN2);
  UB1BPPG_5_3 U5 (O[8], IN1[5], IN2);
  UB1BPPG_6_3 U6 (O[9], IN1[6], IN2);
  UB1BPPG_7_3 U7 (O[10], IN1[7], IN2);
  UB1BPPG_8_3 U8 (O[11], IN1[8], IN2);
  UB1BPPG_9_3 U9 (O[12], IN1[9], IN2);
endmodule

module UBVPPG_9_0_4 (O, IN1, IN2);
  output [13:4] O;
  input [9:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
  UB1BPPG_6_4 U6 (O[10], IN1[6], IN2);
  UB1BPPG_7_4 U7 (O[11], IN1[7], IN2);
  UB1BPPG_8_4 U8 (O[12], IN1[8], IN2);
  UB1BPPG_9_4 U9 (O[13], IN1[9], IN2);
endmodule

module UBVPPG_9_0_5 (O, IN1, IN2);
  output [14:5] O;
  input [9:0] IN1;
  input IN2;
  UB1BPPG_0_5 U0 (O[5], IN1[0], IN2);
  UB1BPPG_1_5 U1 (O[6], IN1[1], IN2);
  UB1BPPG_2_5 U2 (O[7], IN1[2], IN2);
  UB1BPPG_3_5 U3 (O[8], IN1[3], IN2);
  UB1BPPG_4_5 U4 (O[9], IN1[4], IN2);
  UB1BPPG_5_5 U5 (O[10], IN1[5], IN2);
  UB1BPPG_6_5 U6 (O[11], IN1[6], IN2);
  UB1BPPG_7_5 U7 (O[12], IN1[7], IN2);
  UB1BPPG_8_5 U8 (O[13], IN1[8], IN2);
  UB1BPPG_9_5 U9 (O[14], IN1[9], IN2);
endmodule

module UBVPPG_9_0_6 (O, IN1, IN2);
  output [15:6] O;
  input [9:0] IN1;
  input IN2;
  UB1BPPG_0_6 U0 (O[6], IN1[0], IN2);
  UB1BPPG_1_6 U1 (O[7], IN1[1], IN2);
  UB1BPPG_2_6 U2 (O[8], IN1[2], IN2);
  UB1BPPG_3_6 U3 (O[9], IN1[3], IN2);
  UB1BPPG_4_6 U4 (O[10], IN1[4], IN2);
  UB1BPPG_5_6 U5 (O[11], IN1[5], IN2);
  UB1BPPG_6_6 U6 (O[12], IN1[6], IN2);
  UB1BPPG_7_6 U7 (O[13], IN1[7], IN2);
  UB1BPPG_8_6 U8 (O[14], IN1[8], IN2);
  UB1BPPG_9_6 U9 (O[15], IN1[9], IN2);
endmodule

module UBVPPG_9_0_7 (O, IN1, IN2);
  output [16:7] O;
  input [9:0] IN1;
  input IN2;
  UB1BPPG_0_7 U0 (O[7], IN1[0], IN2);
  UB1BPPG_1_7 U1 (O[8], IN1[1], IN2);
  UB1BPPG_2_7 U2 (O[9], IN1[2], IN2);
  UB1BPPG_3_7 U3 (O[10], IN1[3], IN2);
  UB1BPPG_4_7 U4 (O[11], IN1[4], IN2);
  UB1BPPG_5_7 U5 (O[12], IN1[5], IN2);
  UB1BPPG_6_7 U6 (O[13], IN1[6], IN2);
  UB1BPPG_7_7 U7 (O[14], IN1[7], IN2);
  UB1BPPG_8_7 U8 (O[15], IN1[8], IN2);
  UB1BPPG_9_7 U9 (O[16], IN1[9], IN2);
endmodule

module UBVPPG_9_0_8 (O, IN1, IN2);
  output [17:8] O;
  input [9:0] IN1;
  input IN2;
  UB1BPPG_0_8 U0 (O[8], IN1[0], IN2);
  UB1BPPG_1_8 U1 (O[9], IN1[1], IN2);
  UB1BPPG_2_8 U2 (O[10], IN1[2], IN2);
  UB1BPPG_3_8 U3 (O[11], IN1[3], IN2);
  UB1BPPG_4_8 U4 (O[12], IN1[4], IN2);
  UB1BPPG_5_8 U5 (O[13], IN1[5], IN2);
  UB1BPPG_6_8 U6 (O[14], IN1[6], IN2);
  UB1BPPG_7_8 U7 (O[15], IN1[7], IN2);
  UB1BPPG_8_8 U8 (O[16], IN1[8], IN2);
  UB1BPPG_9_8 U9 (O[17], IN1[9], IN2);
endmodule

module UBVPPG_9_0_9 (O, IN1, IN2);
  output [18:9] O;
  input [9:0] IN1;
  input IN2;
  UB1BPPG_0_9 U0 (O[9], IN1[0], IN2);
  UB1BPPG_1_9 U1 (O[10], IN1[1], IN2);
  UB1BPPG_2_9 U2 (O[11], IN1[2], IN2);
  UB1BPPG_3_9 U3 (O[12], IN1[3], IN2);
  UB1BPPG_4_9 U4 (O[13], IN1[4], IN2);
  UB1BPPG_5_9 U5 (O[14], IN1[5], IN2);
  UB1BPPG_6_9 U6 (O[15], IN1[6], IN2);
  UB1BPPG_7_9 U7 (O[16], IN1[7], IN2);
  UB1BPPG_8_9 U8 (O[17], IN1[8], IN2);
  UB1BPPG_9_9 U9 (O[18], IN1[9], IN2);
endmodule

