/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: UBCLA_15_0_63_0

  Operand-1 length: 16
  Operand-2 length: 64
  Two-operand addition algorithm: Carry look-ahead adder
----------------------------------------------------------------------------*/

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_63_16(O);
  output [63:16] O;
  assign O[16] = 0;
  assign O[17] = 0;
  assign O[18] = 0;
  assign O[19] = 0;
  assign O[20] = 0;
  assign O[21] = 0;
  assign O[22] = 0;
  assign O[23] = 0;
  assign O[24] = 0;
  assign O[25] = 0;
  assign O[26] = 0;
  assign O[27] = 0;
  assign O[28] = 0;
  assign O[29] = 0;
  assign O[30] = 0;
  assign O[31] = 0;
  assign O[32] = 0;
  assign O[33] = 0;
  assign O[34] = 0;
  assign O[35] = 0;
  assign O[36] = 0;
  assign O[37] = 0;
  assign O[38] = 0;
  assign O[39] = 0;
  assign O[40] = 0;
  assign O[41] = 0;
  assign O[42] = 0;
  assign O[43] = 0;
  assign O[44] = 0;
  assign O[45] = 0;
  assign O[46] = 0;
  assign O[47] = 0;
  assign O[48] = 0;
  assign O[49] = 0;
  assign O[50] = 0;
  assign O[51] = 0;
  assign O[52] = 0;
  assign O[53] = 0;
  assign O[54] = 0;
  assign O[55] = 0;
  assign O[56] = 0;
  assign O[57] = 0;
  assign O[58] = 0;
  assign O[59] = 0;
  assign O[60] = 0;
  assign O[61] = 0;
  assign O[62] = 0;
  assign O[63] = 0;
endmodule

module GPGenerator(Go, Po, A, B);
  output Go;
  output Po;
  input A;
  input B;
  assign Go = A & B;
  assign Po = A ^ B;
endmodule

module CLAUnit_64(C, G, P, Cin);
  output [64:1] C;
  input Cin;
  input [63:0] G;
  input [63:0] P;
  assign C[1] = G[0] | ( P[0] & Cin );
  assign C[2] = G[1] | ( P[1] & G[0] ) | ( P[1] & P[0] & Cin );
  assign C[3] = G[2] | ( P[2] & G[1] ) | ( P[2] & P[1] & G[0] ) | ( P[2] & P[1] & P[0] & Cin );
  assign C[4] = G[3] | ( P[3] & G[2] ) | ( P[3] & P[2] & G[1] ) | ( P[3] & P[2] & P[1] & G[0] ) | ( P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[5] = G[4] | ( P[4] & G[3] ) | ( P[4] & P[3] & G[2] ) | ( P[4] & P[3] & P[2] & G[1] ) | ( P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[6] = G[5] | ( P[5] & G[4] ) | ( P[5] & P[4] & G[3] ) | ( P[5] & P[4] & P[3] & G[2] ) | ( P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[5] & P[4] & P[3]
 & P[2] & P[1] & P[0] & Cin );
  assign C[7] = G[6] | ( P[6] & G[5] ) | ( P[6] & P[5] & G[4] ) | ( P[6] & P[5] & P[4] & G[3] ) | ( P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[6] & P[5] & P[4]
 & P[3] & P[2] & P[1] & G[0] ) | ( P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[8] = G[7] | ( P[7] & G[6] ) | ( P[7] & P[6] & G[5] ) | ( P[7] & P[6] & P[5] & G[4] ) | ( P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[7] & P[6] & P[5]
 & P[4] & P[3] & P[2] & G[1] ) | ( P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[9] = G[8] | ( P[8] & G[7] ) | ( P[8] & P[7] & G[6] ) | ( P[8] & P[7] & P[6] & G[5] ) | ( P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & G[2] ) | ( P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[8] & P[7] & P[6] & P[5] & P[4] & P[3]
 & P[2] & P[1] & P[0] & Cin );
  assign C[10] = G[9] | ( P[9] & G[8] ) | ( P[9] & P[8] & G[7] ) | ( P[9] & P[8] & P[7] & G[6] ) | ( P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & G[3] ) | ( P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & P[1] & G[0] ) | ( P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[11] = G[10] | ( P[10] & G[9] ) | ( P[10] & P[9] & G[8] ) | ( P[10] & P[9] & P[8] & G[7] ) | ( P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] &
 Cin );
  assign C[12] = G[11] | ( P[11] & G[10] ) | ( P[11] & P[10] & G[9] ) | ( P[11] & P[10] & P[9] & G[8] ) | ( P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[11]
 & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[11] & P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3]
 & P[2] & P[1] & G[0] ) | ( P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[13] = G[12] | ( P[12] & G[11] ) | ( P[12] & P[11] & G[10] ) | ( P[12] & P[11] & P[10] & G[9] ) | ( P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & G[1] ) | ( P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2]
 & P[1] & P[0] & Cin );
  assign C[14] = G[13] | ( P[13] & G[12] ) | ( P[13] & P[12] & G[11] ) | ( P[13] & P[12] & P[11] & G[10] ) | ( P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) |
 ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[13] &
 P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] &
 P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[15] = G[14] | ( P[14] & G[13] ) | ( P[14] & P[13] & G[12] ) | ( P[14] & P[13] & P[12] & G[11] ) | ( P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & G[9] )
 | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] &
 P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[16] = G[15] | ( P[15] & G[14] ) | ( P[15] & P[14] & G[13] ) | ( P[15] & P[14] & P[13] & G[12] ) | ( P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & G[10] )
 | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | (
 P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[15] & P[14] & P[13] &
 P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] &
 P[1] & P[0] & Cin );
  assign C[17] = G[16] | ( P[16] & G[15] ) | ( P[16] & P[15] & G[14] ) | ( P[16] & P[15] & P[14] & G[13] ) | ( P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & G[11] )
 | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] )
 | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[16] & P[15]
 & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & P[1] & G[0] ) | ( P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[18] = G[17] | ( P[17] & G[16] ) | ( P[17] & P[16] & G[15] ) | ( P[17] & P[16] & P[15] & G[14] ) | ( P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & G[12] )
 | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9]
 ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[17] & P[16] &
 P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[19] = G[18] | ( P[18] & G[17] ) | ( P[18] & P[17] & G[16] ) | ( P[18] & P[17] & P[16] & G[15] ) | ( P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & G[13] )
 | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10]
 ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4]
 ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | (
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] &
 P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[20] = G[19] | ( P[19] & G[18] ) | ( P[19] & P[18] & G[17] ) | ( P[19] & P[18] & P[17] & G[16] ) | ( P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & G[14] )
 | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11]
 ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5]
 ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) |
 ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] &
 P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[21] = G[20] | ( P[20] & G[19] ) | ( P[20] & P[19] & G[18] ) | ( P[20] & P[19] & P[18] & G[17] ) | ( P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & G[15] )
 | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12]
 ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6]
 ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] )
 | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8]
 & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2]
 & P[1] & P[0] & Cin );
  assign C[22] = G[21] | ( P[21] & G[20] ) | ( P[21] & P[20] & G[19] ) | ( P[21] & P[20] & P[19] & G[18] ) | ( P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & G[16] )
 | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13]
 ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[21] & P[20] & P[19]
 & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] &
 P[8] & G[7] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & G[4] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] &
 P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2]
 & P[1] & P[0] & Cin );
  assign C[23] = G[22] | ( P[22] & G[21] ) | ( P[22] & P[21] & G[20] ) | ( P[22] & P[21] & P[20] & G[19] ) | ( P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & G[17] )
 | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14]
 ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & G[8] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & G[5] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8]
 & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] &
 P[3] & P[2] & P[1] & G[0] ) | ( P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0]
 & Cin );
  assign C[24] = G[23] | ( P[23] & G[22] ) | ( P[23] & P[22] & G[21] ) | ( P[23] & P[22] & P[21] & G[20] ) | ( P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & G[18] )
 | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15]
 ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & G[9] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] &
 P[8] & P[7] & G[6] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] &
 P[4] & P[3] & P[2] & G[1] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1]
 & G[0] ) | ( P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[25] = G[24] | ( P[24] & G[23] ) | ( P[24] & P[23] & G[22] ) | ( P[24] & P[23] & P[22] & G[21] ) | ( P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & G[19] )
 | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16]
 ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & G[10] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] &
 P[10] & P[9] & P[8] & G[7] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8]
 & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5]
 & P[4] & P[3] & P[2] & G[1] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3]
 & P[2] & P[1] & G[0] ) | ( P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2]
 & P[1] & P[0] & Cin );
  assign C[26] = G[25] | ( P[25] & G[24] ) | ( P[25] & P[24] & G[23] ) | ( P[25] & P[24] & P[23] & G[22] ) | ( P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & G[20] )
 | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17]
 ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & G[11] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & G[8] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5]
 & P[4] & P[3] & P[2] & G[1] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & P[1] & G[0] ) | ( P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[27] = G[26] | ( P[26] & G[25] ) | ( P[26] & P[25] & G[24] ) | ( P[26] & P[25] & P[24] & G[23] ) | ( P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & G[21] )
 | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18]
 ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[26] & P[25] &
 P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & G[12] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & G[9] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] &
 P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[28] = G[27] | ( P[27] & G[26] ) | ( P[27] & P[26] & G[25] ) | ( P[27] & P[26] & P[25] & G[24] ) | ( P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & G[22] )
 | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19]
 ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[27] & P[26] &
 P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & G[13] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & G[10] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] &
 P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[29] = G[28] | ( P[28] & G[27] ) | ( P[28] & P[27] & G[26] ) | ( P[28] & P[27] & P[26] & G[25] ) | ( P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & G[23] )
 | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20]
 ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & G[14] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & P[13] & P[12] & G[11] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19]
 & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[30] = G[29] | ( P[29] & G[28] ) | ( P[29] & P[28] & G[27] ) | ( P[29] & P[28] & P[27] & G[26] ) | ( P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & G[24] )
 | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21]
 ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[29] & P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & G[15] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & G[12] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19]
 & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[31] = G[30] | ( P[30] & G[29] ) | ( P[30] & P[29] & G[28] ) | ( P[30] & P[29] & P[28] & G[27] ) | ( P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & G[25] )
 | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22]
 ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & G[16] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] &
 P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & G[13] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[30] &
 P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[32] = G[31] | ( P[31] & G[30] ) | ( P[31] & P[30] & G[29] ) | ( P[31] & P[30] & P[29] & G[28] ) | ( P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & G[26] )
 | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23]
 ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[31] & P[30] &
 P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19]
 & P[18] & G[17] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] &
 P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & G[14] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[31] &
 P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19]
 & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] &
 P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] )
 | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] &
 P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[33] = G[32] | ( P[32] & G[31] ) | ( P[32] & P[31] & G[30] ) | ( P[32] & P[31] & P[30] & G[29] ) | ( P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & G[27] )
 | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24]
 ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[32] & P[31] &
 P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & G[18] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19]
 & P[18] & P[17] & P[16] & G[15] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[32] &
 P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3]
 & G[2] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9]
 & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[34] = G[33] | ( P[33] & G[32] ) | ( P[33] & P[32] & G[31] ) | ( P[33] & P[32] & P[31] & G[30] ) | ( P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & G[28] )
 | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25]
 ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[33] & P[32] &
 P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & G[19] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & G[16] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[33] &
 P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19]
 & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19]
 & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5]
 & P[4] & G[3] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[35] = G[34] | ( P[34] & G[33] ) | ( P[34] & P[33] & G[32] ) | ( P[34] & P[33] & P[32] & G[31] ) | ( P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & G[29] )
 | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26]
 ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[34] & P[33] &
 P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & G[20] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & G[17] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[34] &
 P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19]
 & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19]
 & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & G[4] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19]
 & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] &
 P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[36] = G[35] | ( P[35] & G[34] ) | ( P[35] & P[34] & G[33] ) | ( P[35] & P[34] & P[33] & G[32] ) | ( P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & G[30] )
 | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27]
 ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[35] & P[34] &
 P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & G[21] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] &
 P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & G[18] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[35] &
 P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[35] &
 P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9]
 & P[8] & P[7] & P[6] & G[5] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] )
 | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[37] = G[36] | ( P[36] & G[35] ) | ( P[36] & P[35] & G[34] ) | ( P[36] & P[35] & P[34] & G[33] ) | ( P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & G[31] )
 | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28]
 ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[36] & P[35] &
 P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & G[22] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] &
 P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & G[19] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[36] &
 P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] &
 P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & G[3] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[38] = G[37] | ( P[37] & G[36] ) | ( P[37] & P[36] & G[35] ) | ( P[37] & P[36] & P[35] & G[34] ) | ( P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & G[32] )
 | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29]
 ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[37] & P[36] &
 P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & G[23] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] &
 P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & G[20] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[37] &
 P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] &
 P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] &
 P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & G[4] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] &
 P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[39] = G[38] | ( P[38] & G[37] ) | ( P[38] & P[37] & G[36] ) | ( P[38] & P[37] & P[36] & G[35] ) | ( P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & G[33] )
 | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30]
 ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[38] & P[37] &
 P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & G[24] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] &
 P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & G[21] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[38] &
 P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] &
 P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] &
 P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & G[5] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] &
 P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[40] = G[39] | ( P[39] & G[38] ) | ( P[39] & P[38] & G[37] ) | ( P[39] & P[38] & P[37] & G[36] ) | ( P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & G[34] )
 | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31]
 ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[39] & P[38] &
 P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & G[25] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] &
 P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & G[22] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[39] &
 P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] &
 P[9] & P[8] & P[7] & G[6] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] &
 P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] &
 P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] &
 P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[41] = G[40] | ( P[40] & G[39] ) | ( P[40] & P[39] & G[38] ) | ( P[40] & P[39] & P[38] & G[37] ) | ( P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & G[35] )
 | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32]
 ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[40] & P[39] &
 P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & G[26] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] &
 P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & G[23] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[40] &
 P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] &
 P[10] & P[9] & P[8] & G[7] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[40] &
 P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] &
 P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] &
 P[2] & P[1] & P[0] & Cin );
  assign C[42] = G[41] | ( P[41] & G[40] ) | ( P[41] & P[40] & G[39] ) | ( P[41] & P[40] & P[39] & G[38] ) | ( P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & G[36] )
 | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33]
 ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[41] & P[40] &
 P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & G[27] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] &
 P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & G[24] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[41] &
 P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] &
 P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] &
 P[11] & P[10] & P[9] & G[8] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] &
 P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] &
 P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] &
 P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5]
 & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[43] = G[42] | ( P[42] & G[41] ) | ( P[42] & P[41] & G[40] ) | ( P[42] & P[41] & P[40] & G[39] ) | ( P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & G[37] )
 | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34]
 ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[42] & P[41] &
 P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & G[28] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] &
 P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & G[25] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[42] &
 P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] &
 P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] &
 P[12] & P[11] & P[10] & G[9] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) |
 ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[42] &
 P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]
 ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[44] = G[43] | ( P[43] & G[42] ) | ( P[43] & P[42] & G[41] ) | ( P[43] & P[42] & P[41] & G[40] ) | ( P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & G[38] )
 | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35]
 ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[43] & P[42] &
 P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & G[29] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] &
 P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & G[26] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[43] &
 P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & G[10] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) |
 ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] &
 P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5]
 & G[4] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] &
 P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] &
 P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[45] = G[44] | ( P[44] & G[43] ) | ( P[44] & P[43] & G[42] ) | ( P[44] & P[43] & P[42] & G[41] ) | ( P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & G[39] )
 | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36]
 ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[44] & P[43] &
 P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & G[30] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] &
 P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & G[27] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[44] &
 P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & G[11] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] )
 | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) |
 ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & G[5] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] &
 P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] )
 | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] &
 P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] &
 P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[46] = G[45] | ( P[45] & G[44] ) | ( P[45] & P[44] & G[43] ) | ( P[45] & P[44] & P[43] & G[42] ) | ( P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & G[40] )
 | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37]
 ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[45] & P[44] &
 P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & G[31] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] &
 P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & G[28] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[45] &
 P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] &
 P[15] & P[14] & P[13] & G[12] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] )
 | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) |
 ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] &
 P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9]
 & P[8] & P[7] & G[6] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] &
 P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & G[3] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] &
 P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3]
 & P[2] & P[1] & P[0] & Cin );
  assign C[47] = G[46] | ( P[46] & G[45] ) | ( P[46] & P[45] & G[44] ) | ( P[46] & P[45] & P[44] & G[43] ) | ( P[46] & P[45] & P[44] & P[43] & G[42] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & G[41] )
 | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38]
 ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[46] & P[45] &
 P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & G[32] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] &
 P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & G[29] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[46] &
 P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] &
 P[16] & P[15] & P[14] & G[13] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] )
 | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] )
 | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] &
 P[10] & P[9] & P[8] & G[7] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] &
 P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] &
 P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & G[4] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] &
 P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] &
 P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5]
 & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0]
 & Cin );
  assign C[48] = G[47] | ( P[47] & G[46] ) | ( P[47] & P[46] & G[45] ) | ( P[47] & P[46] & P[45] & G[44] ) | ( P[47] & P[46] & P[45] & P[44] & G[43] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & G[42] )
 | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39]
 ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[47] & P[46] &
 P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & G[33] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] &
 P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & G[30] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[47] &
 P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & G[14] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] )
 | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] )
 | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23]
 & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] &
 P[11] & P[10] & P[9] & G[8] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] &
 P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17]
 & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] &
 P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8]
 & P[7] & P[6] & G[5] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] &
 P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] &
 P[1] & G[0] ) | ( P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] &
 P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[49] = G[48] | ( P[48] & G[47] ) | ( P[48] & P[47] & G[46] ) | ( P[48] & P[47] & P[46] & G[45] ) | ( P[48] & P[47] & P[46] & P[45] & G[44] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & G[43] )
 | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & G[42] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40]
 ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[48] & P[47] &
 P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & G[34] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] &
 P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & G[31] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[48] &
 P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & G[15] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] )
 | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] )
 | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] &
 P[12] & P[11] & P[10] & G[9] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] &
 P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & G[6] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] &
 P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5]
 & P[4] & P[3] & P[2] & G[1] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1]
 & G[0] ) | ( P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[50] = G[49] | ( P[49] & G[48] ) | ( P[49] & P[48] & G[47] ) | ( P[49] & P[48] & P[47] & G[46] ) | ( P[49] & P[48] & P[47] & P[46] & G[45] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & G[44] )
 | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & G[43] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & G[42] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41]
 ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[49] & P[48] &
 P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & G[35] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] &
 P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & G[32] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[49] &
 P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & G[16] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] )
 | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] )
 | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & G[10] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] &
 P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & P[9] & P[8] & G[7] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[49] & P[48] &
 P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] &
 P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] &
 P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & G[2] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] &
 P[2] & G[1] ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]
 ) | ( P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[51] = G[50] | ( P[50] & G[49] ) | ( P[50] & P[49] & G[48] ) | ( P[50] & P[49] & P[48] & G[47] ) | ( P[50] & P[49] & P[48] & P[47] & G[46] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & G[45] )
 | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & G[44] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & G[43] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & G[42]
 ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[50] & P[49] &
 P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & G[36] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] &
 P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & G[33] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[50] &
 P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] &
 P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & G[17] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] )
 | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] )
 | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & G[11] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] &
 P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] &
 P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[50] &
 P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] &
 P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] &
 P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13]
 & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] &
 P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5]
 & P[4] & P[3] & G[2] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3]
 & P[2] & G[1] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] &
 P[1] & G[0] ) | ( P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1]
 & P[0] & Cin );
  assign C[52] = G[51] | ( P[51] & G[50] ) | ( P[51] & P[50] & G[49] ) | ( P[51] & P[50] & P[49] & G[48] ) | ( P[51] & P[50] & P[49] & P[48] & G[47] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & G[46] )
 | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & G[45] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & G[44] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & G[43]
 ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & G[42] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[51] & P[50] &
 P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & G[37] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] &
 P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & G[34] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[51] &
 P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] &
 P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & G[18] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] )
 | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] )
 | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] &
 P[15] & P[14] & P[13] & G[12] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] &
 P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] &
 P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] &
 P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] &
 P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & G[3] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] &
 P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5]
 & P[4] & P[3] & G[2] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & G[1] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4]
 & P[3] & P[2] & P[1] & G[0] ) | ( P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] &
 P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5]
 & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[53] = G[52] | ( P[52] & G[51] ) | ( P[52] & P[51] & G[50] ) | ( P[52] & P[51] & P[50] & G[49] ) | ( P[52] & P[51] & P[50] & P[49] & G[48] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & G[47] )
 | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & G[46] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & G[45] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & G[44]
 ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & G[43] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & G[42] ) | ( P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[52] & P[51] &
 P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & G[38] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] &
 P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & G[35] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[52] &
 P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & G[19] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] )
 | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] )
 | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28]
 & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] &
 P[16] & P[15] & P[14] & G[13] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] &
 P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] &
 P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] &
 P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] &
 P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & G[3] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] &
 P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & G[2] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] &
 P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] &
 P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] &
 P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[54] = G[53] | ( P[53] & G[52] ) | ( P[53] & P[52] & G[51] ) | ( P[53] & P[52] & P[51] & G[50] ) | ( P[53] & P[52] & P[51] & P[50] & G[49] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & G[48] )
 | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & G[47] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & G[46] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & G[45]
 ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & G[44] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & G[43] ) | ( P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & G[42] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[53] & P[52] &
 P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & G[39] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] &
 P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & G[36] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[53] &
 P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] &
 P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & G[20] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] )
 | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] )
 | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & G[14] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] &
 P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] &
 P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] &
 P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] &
 P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] &
 P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] &
 P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] &
 P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] &
 P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] &
 P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[55] = G[54] | ( P[54] & G[53] ) | ( P[54] & P[53] & G[52] ) | ( P[54] & P[53] & P[52] & G[51] ) | ( P[54] & P[53] & P[52] & P[51] & G[50] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & G[49] )
 | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & G[48] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & G[47] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & G[46]
 ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & G[45] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & G[44] ) | ( P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & G[43] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & G[42] ) | ( P[54] & P[53] &
 P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & G[40] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] &
 P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & G[37] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[54] &
 P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] &
 P[24] & P[23] & P[22] & G[21] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] )
 | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] )
 | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & G[15] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] &
 P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] &
 P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] &
 P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] &
 P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] &
 P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] &
 P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] &
 P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] &
 P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] &
 P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20]
 & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[56] = G[55] | ( P[55] & G[54] ) | ( P[55] & P[54] & G[53] ) | ( P[55] & P[54] & P[53] & G[52] ) | ( P[55] & P[54] & P[53] & P[52] & G[51] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & G[50] )
 | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & G[49] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & G[48] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & G[47]
 ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & G[46] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & G[45] ) | ( P[55] & P[54] & P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & G[44] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & G[43] ) | ( P[55] & P[54] &
 P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & G[42] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & G[41] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] &
 P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & G[38] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[55] &
 P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[55]
 & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] &
 P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] &
 P[25] & P[24] & P[23] & G[22] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] )
 | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] )
 | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & G[16] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] &
 P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[55]
 & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] &
 P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] &
 P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] &
 P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] &
 P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] &
 P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] &
 P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[55] & P[54] & P[53] &
 P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27]
 & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] &
 P[0] & Cin );
  assign C[57] = G[56] | ( P[56] & G[55] ) | ( P[56] & P[55] & G[54] ) | ( P[56] & P[55] & P[54] & G[53] ) | ( P[56] & P[55] & P[54] & P[53] & G[52] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & G[51] )
 | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & G[50] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & G[49] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & G[48]
 ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & G[47] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & G[46] ) | ( P[56] & P[55] & P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & G[45] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & G[44] ) | ( P[56] & P[55] &
 P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & G[43] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & G[42] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] &
 P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & G[39] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[56] &
 P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[56]
 & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] &
 P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[56] & P[55] & P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & G[23] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] )
 | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] )
 | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]
 & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & G[17] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[56] & P[55] & P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[56]
 & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] &
 P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] &
 P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] &
 P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] &
 P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] &
 P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] &
 P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[56] & P[55]
 & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] &
 P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] &
 P[3] & P[2] & P[1] & G[0] ) | ( P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] &
 P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[58] = G[57] | ( P[57] & G[56] ) | ( P[57] & P[56] & G[55] ) | ( P[57] & P[56] & P[55] & G[54] ) | ( P[57] & P[56] & P[55] & P[54] & G[53] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & G[52] )
 | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & G[51] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & G[50] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & G[49]
 ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & G[48] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & G[47] ) | ( P[57] & P[56] & P[55]
 & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & G[46] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & G[45] ) | ( P[57] & P[56] &
 P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & G[44] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & G[43] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & G[42] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] &
 P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & G[40] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[57] &
 P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[57]
 & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] &
 P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[57] & P[56] & P[55] & P[54] & P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] &
 P[27] & P[26] & P[25] & G[24] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] )
 | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] )
 | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33]
 & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & G[18] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[57] & P[56] & P[55] & P[54] & P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[57]
 & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] &
 P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] &
 P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] &
 P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] &
 P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[57]
 & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] &
 P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] &
 P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[59] = G[58] | ( P[58] & G[57] ) | ( P[58] & P[57] & G[56] ) | ( P[58] & P[57] & P[56] & G[55] ) | ( P[58] & P[57] & P[56] & P[55] & G[54] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & G[53] )
 | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & G[52] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & G[51] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & G[50]
 ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & G[49] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & G[48] ) | ( P[58] & P[57] & P[56]
 & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & G[47] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & G[46] ) | ( P[58] & P[57] &
 P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & G[45] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & G[44] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & G[43] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] &
 P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & G[42] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & G[41] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[58] &
 P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[58]
 & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] &
 P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[58] & P[57] & P[56] & P[55] & P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] &
 P[28] & P[27] & P[26] & G[25] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] )
 | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] )
 | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & G[19] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[58] & P[57] & P[56] & P[55] & P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[58]
 & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] &
 P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] &
 P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] &
 P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[58] & P[57] & P[56] & P[55] & P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] )
 | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34]
 & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] &
 P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[58] & P[57] & P[56] & P[55] &
 P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3]
 & P[2] & P[1] & P[0] & Cin );
  assign C[60] = G[59] | ( P[59] & G[58] ) | ( P[59] & P[58] & G[57] ) | ( P[59] & P[58] & P[57] & G[56] ) | ( P[59] & P[58] & P[57] & P[56] & G[55] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & G[54] )
 | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & G[53] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & G[52] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & G[51]
 ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & G[50] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & G[49] ) | ( P[59] & P[58] & P[57]
 & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & G[48] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & G[47] ) | ( P[59] & P[58] &
 P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & G[46] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & G[45] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & G[44] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] &
 P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & G[43] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & G[42] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[59] &
 P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[59]
 & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] &
 P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[59] & P[58] & P[57] & P[56] & P[55]
 & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] &
 P[29] & P[28] & P[27] & G[26] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] )
 | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] )
 | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35]
 & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & G[20] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[59] & P[58] & P[57] & P[56] & P[55]
 & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] &
 P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[59]
 & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] &
 P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] &
 P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] &
 P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21]
 & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[59] & P[58] & P[57] & P[56]
 & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] &
 P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5]
 & G[4] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] &
 P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] &
 P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[59] & P[58] & P[57]
 & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] &
 P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6]
 & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[61] = G[60] | ( P[60] & G[59] ) | ( P[60] & P[59] & G[58] ) | ( P[60] & P[59] & P[58] & G[57] ) | ( P[60] & P[59] & P[58] & P[57] & G[56] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & G[55] )
 | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & G[54] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & G[53] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & G[52]
 ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & G[51] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & G[50] ) | ( P[60] & P[59] & P[58]
 & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & G[49] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & G[48] ) | ( P[60] & P[59] &
 P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & G[47] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & G[46] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & G[45] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] &
 P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & G[44] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & G[43] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & G[42] ) | ( P[60] &
 P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55]
 & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55]
 & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[60]
 & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] &
 P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[60] & P[59] & P[58] & P[57] & P[56]
 & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] &
 P[30] & P[29] & P[28] & G[27] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] )
 | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] )
 | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] &
 P[24] & P[23] & P[22] & G[21] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[60] & P[59] & P[58] & P[57] & P[56]
 & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] &
 P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[60]
 & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] &
 P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55]
 & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] &
 P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] &
 P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] &
 P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25]
 & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[60] & P[59] & P[58]
 & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] &
 P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & G[5] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] &
 P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] &
 P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[60] & P[59]
 & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] &
 P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8]
 & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] &
 P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] &
 P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26]
 & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin
 );
  assign C[62] = G[61] | ( P[61] & G[60] ) | ( P[61] & P[60] & G[59] ) | ( P[61] & P[60] & P[59] & G[58] ) | ( P[61] & P[60] & P[59] & P[58] & G[57] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & G[56] )
 | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & G[55] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & G[54] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & G[53]
 ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & G[52] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & G[51] ) | ( P[61] & P[60] & P[59]
 & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & G[50] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & G[49] ) | ( P[61] & P[60] &
 P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & G[48] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & G[47] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & G[46] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] &
 P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & G[45] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & G[44] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & G[43] ) | ( P[61] &
 P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & G[42] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56]
 & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56]
 & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[61]
 & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] &
 P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[61] & P[60] & P[59] & P[58] & P[57]
 & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] &
 P[31] & P[30] & P[29] & G[28] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] )
 | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] )
 | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37]
 & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] &
 P[25] & P[24] & P[23] & G[22] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41]
 & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[61] & P[60] & P[59] & P[58] & P[57]
 & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] &
 P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[61]
 & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] &
 P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56]
 & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] &
 P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] &
 P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30]
 & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[61] & P[60]
 & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] &
 P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9]
 & P[8] & P[7] & G[6] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40]
 & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] &
 P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46]
 & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] &
 P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[61]
 & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] &
 P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10]
 & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] &
 P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] &
 P[2] & P[1] & G[0] ) | ( P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] &
 P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14]
 & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
  assign C[63] = G[62] | ( P[62] & G[61] ) | ( P[62] & P[61] & G[60] ) | ( P[62] & P[61] & P[60] & G[59] ) | ( P[62] & P[61] & P[60] & P[59] & G[58] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & G[57] )
 | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & G[56] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & G[55] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & G[54]
 ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & G[53] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & G[52] ) | ( P[62] & P[61] & P[60]
 & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & G[51] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & G[50] ) | ( P[62] & P[61] &
 P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & G[49] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & G[48] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & G[47] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] &
 P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & G[46] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & G[45] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & G[44] ) | ( P[62] &
 P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & G[43] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57]
 & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & G[42] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57]
 & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[62]
 & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] &
 P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & G[30] ) | ( P[62] & P[61] & P[60] & P[59] & P[58]
 & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] &
 P[32] & P[31] & P[30] & G[29] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] )
 | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] )
 | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38]
 & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & G[24] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & G[23] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[62] & P[61] & P[60] & P[59] & P[58]
 & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] &
 P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] &
 P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[62]
 & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] &
 P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57]
 & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] &
 P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] &
 P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47]
 & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] &
 P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] &
 P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] &
 P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57]
 & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] &
 P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8] ) | ( P[62] &
 P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36]
 & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] &
 P[10] & P[9] & P[8] & G[7] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] &
 P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16]
 & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] &
 P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22]
 & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] &
 P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29]
 & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[62]
 & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] &
 P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11]
 & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45]
 & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] &
 P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55]
 & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] &
 P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] &
 P[3] & P[2] & G[1] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] &
 P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15]
 & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0] ) | ( P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52]
 & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] &
 P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0]
 & Cin );
  assign C[64] = G[63] | ( P[63] & G[62] ) | ( P[63] & P[62] & G[61] ) | ( P[63] & P[62] & P[61] & G[60] ) | ( P[63] & P[62] & P[61] & P[60] & G[59] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & G[58] )
 | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & G[57] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & G[56] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & G[55]
 ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & G[54] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & G[53] ) | ( P[63] & P[62] & P[61]
 & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & G[52] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & G[51] ) | ( P[63] & P[62] &
 P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & G[50] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & G[49] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & G[48] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] &
 P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & G[47] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50]
 & P[49] & P[48] & P[47] & G[46] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & G[45] ) | ( P[63] &
 P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & G[44] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58]
 & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & G[43] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & G[42] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & G[41] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & G[40] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & G[39] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & G[38] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & G[37] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & G[36] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & G[35] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58]
 & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & G[34] ) | ( P[63]
 & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] &
 P[37] & P[36] & P[35] & P[34] & G[33] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & G[32] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & G[31] ) | ( P[63] & P[62] & P[61] & P[60] & P[59]
 & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] &
 P[33] & P[32] & P[31] & G[30] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & G[29] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & G[28] )
 | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & G[27] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & G[26] )
 | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & G[25] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53]
 & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] &
 P[27] & P[26] & P[25] & G[24] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & G[23] ) | ( P[63] & P[62] & P[61] & P[60] & P[59]
 & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] &
 P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & G[22] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] &
 P[25] & P[24] & P[23] & P[22] & G[21] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44]
 & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & G[20] ) | ( P[63]
 & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] &
 P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & G[19] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58]
 & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] &
 P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & G[18] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & G[17] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] &
 P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & G[16] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & G[15] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & G[14] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & G[13] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49]
 & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] &
 P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & G[12] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51]
 & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] &
 P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & G[11] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54]
 & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] &
 P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & G[10] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58]
 & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] &
 P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9] ) | ( P[63]
 & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] &
 P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12]
 & P[11] & P[10] & P[9] & G[8] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43]
 & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] &
 P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] &
 P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24]
 & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] &
 P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31]
 & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5]
 ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39]
 & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] &
 P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48]
 & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] &
 P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58]
 & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] &
 P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7]
 & P[6] & P[5] & P[4] & P[3] & G[2] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] &
 P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18]
 & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55]
 & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] &
 P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] & P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] &
 P[3] & P[2] & P[1] & G[0] ) | ( P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42]
 & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32] & P[31] & P[30] & P[29] & P[28] & P[27] & P[26] & P[25] & P[24] & P[23] & P[22] & P[21] & P[20] & P[19] & P[18] & P[17] &
 P[16] & P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin );
endmodule

module UBPriCLA_63_0(S, X, Y, Cin);
  output [64:0] S;
  input Cin;
  input [63:0] X;
  input [63:0] Y;
  wire [64:1] C;
  wire [63:0] G;
  wire [63:0] P;
  assign S[0] = Cin ^ P[0];
  assign S[1] = C[1] ^ P[1];
  assign S[2] = C[2] ^ P[2];
  assign S[3] = C[3] ^ P[3];
  assign S[4] = C[4] ^ P[4];
  assign S[5] = C[5] ^ P[5];
  assign S[6] = C[6] ^ P[6];
  assign S[7] = C[7] ^ P[7];
  assign S[8] = C[8] ^ P[8];
  assign S[9] = C[9] ^ P[9];
  assign S[10] = C[10] ^ P[10];
  assign S[11] = C[11] ^ P[11];
  assign S[12] = C[12] ^ P[12];
  assign S[13] = C[13] ^ P[13];
  assign S[14] = C[14] ^ P[14];
  assign S[15] = C[15] ^ P[15];
  assign S[16] = C[16] ^ P[16];
  assign S[17] = C[17] ^ P[17];
  assign S[18] = C[18] ^ P[18];
  assign S[19] = C[19] ^ P[19];
  assign S[20] = C[20] ^ P[20];
  assign S[21] = C[21] ^ P[21];
  assign S[22] = C[22] ^ P[22];
  assign S[23] = C[23] ^ P[23];
  assign S[24] = C[24] ^ P[24];
  assign S[25] = C[25] ^ P[25];
  assign S[26] = C[26] ^ P[26];
  assign S[27] = C[27] ^ P[27];
  assign S[28] = C[28] ^ P[28];
  assign S[29] = C[29] ^ P[29];
  assign S[30] = C[30] ^ P[30];
  assign S[31] = C[31] ^ P[31];
  assign S[32] = C[32] ^ P[32];
  assign S[33] = C[33] ^ P[33];
  assign S[34] = C[34] ^ P[34];
  assign S[35] = C[35] ^ P[35];
  assign S[36] = C[36] ^ P[36];
  assign S[37] = C[37] ^ P[37];
  assign S[38] = C[38] ^ P[38];
  assign S[39] = C[39] ^ P[39];
  assign S[40] = C[40] ^ P[40];
  assign S[41] = C[41] ^ P[41];
  assign S[42] = C[42] ^ P[42];
  assign S[43] = C[43] ^ P[43];
  assign S[44] = C[44] ^ P[44];
  assign S[45] = C[45] ^ P[45];
  assign S[46] = C[46] ^ P[46];
  assign S[47] = C[47] ^ P[47];
  assign S[48] = C[48] ^ P[48];
  assign S[49] = C[49] ^ P[49];
  assign S[50] = C[50] ^ P[50];
  assign S[51] = C[51] ^ P[51];
  assign S[52] = C[52] ^ P[52];
  assign S[53] = C[53] ^ P[53];
  assign S[54] = C[54] ^ P[54];
  assign S[55] = C[55] ^ P[55];
  assign S[56] = C[56] ^ P[56];
  assign S[57] = C[57] ^ P[57];
  assign S[58] = C[58] ^ P[58];
  assign S[59] = C[59] ^ P[59];
  assign S[60] = C[60] ^ P[60];
  assign S[61] = C[61] ^ P[61];
  assign S[62] = C[62] ^ P[62];
  assign S[63] = C[63] ^ P[63];
  assign S[64] = C[64];
  GPGenerator U0 (G[0], P[0], X[0], Y[0]);
  GPGenerator U1 (G[1], P[1], X[1], Y[1]);
  GPGenerator U2 (G[2], P[2], X[2], Y[2]);
  GPGenerator U3 (G[3], P[3], X[3], Y[3]);
  GPGenerator U4 (G[4], P[4], X[4], Y[4]);
  GPGenerator U5 (G[5], P[5], X[5], Y[5]);
  GPGenerator U6 (G[6], P[6], X[6], Y[6]);
  GPGenerator U7 (G[7], P[7], X[7], Y[7]);
  GPGenerator U8 (G[8], P[8], X[8], Y[8]);
  GPGenerator U9 (G[9], P[9], X[9], Y[9]);
  GPGenerator U10 (G[10], P[10], X[10], Y[10]);
  GPGenerator U11 (G[11], P[11], X[11], Y[11]);
  GPGenerator U12 (G[12], P[12], X[12], Y[12]);
  GPGenerator U13 (G[13], P[13], X[13], Y[13]);
  GPGenerator U14 (G[14], P[14], X[14], Y[14]);
  GPGenerator U15 (G[15], P[15], X[15], Y[15]);
  GPGenerator U16 (G[16], P[16], X[16], Y[16]);
  GPGenerator U17 (G[17], P[17], X[17], Y[17]);
  GPGenerator U18 (G[18], P[18], X[18], Y[18]);
  GPGenerator U19 (G[19], P[19], X[19], Y[19]);
  GPGenerator U20 (G[20], P[20], X[20], Y[20]);
  GPGenerator U21 (G[21], P[21], X[21], Y[21]);
  GPGenerator U22 (G[22], P[22], X[22], Y[22]);
  GPGenerator U23 (G[23], P[23], X[23], Y[23]);
  GPGenerator U24 (G[24], P[24], X[24], Y[24]);
  GPGenerator U25 (G[25], P[25], X[25], Y[25]);
  GPGenerator U26 (G[26], P[26], X[26], Y[26]);
  GPGenerator U27 (G[27], P[27], X[27], Y[27]);
  GPGenerator U28 (G[28], P[28], X[28], Y[28]);
  GPGenerator U29 (G[29], P[29], X[29], Y[29]);
  GPGenerator U30 (G[30], P[30], X[30], Y[30]);
  GPGenerator U31 (G[31], P[31], X[31], Y[31]);
  GPGenerator U32 (G[32], P[32], X[32], Y[32]);
  GPGenerator U33 (G[33], P[33], X[33], Y[33]);
  GPGenerator U34 (G[34], P[34], X[34], Y[34]);
  GPGenerator U35 (G[35], P[35], X[35], Y[35]);
  GPGenerator U36 (G[36], P[36], X[36], Y[36]);
  GPGenerator U37 (G[37], P[37], X[37], Y[37]);
  GPGenerator U38 (G[38], P[38], X[38], Y[38]);
  GPGenerator U39 (G[39], P[39], X[39], Y[39]);
  GPGenerator U40 (G[40], P[40], X[40], Y[40]);
  GPGenerator U41 (G[41], P[41], X[41], Y[41]);
  GPGenerator U42 (G[42], P[42], X[42], Y[42]);
  GPGenerator U43 (G[43], P[43], X[43], Y[43]);
  GPGenerator U44 (G[44], P[44], X[44], Y[44]);
  GPGenerator U45 (G[45], P[45], X[45], Y[45]);
  GPGenerator U46 (G[46], P[46], X[46], Y[46]);
  GPGenerator U47 (G[47], P[47], X[47], Y[47]);
  GPGenerator U48 (G[48], P[48], X[48], Y[48]);
  GPGenerator U49 (G[49], P[49], X[49], Y[49]);
  GPGenerator U50 (G[50], P[50], X[50], Y[50]);
  GPGenerator U51 (G[51], P[51], X[51], Y[51]);
  GPGenerator U52 (G[52], P[52], X[52], Y[52]);
  GPGenerator U53 (G[53], P[53], X[53], Y[53]);
  GPGenerator U54 (G[54], P[54], X[54], Y[54]);
  GPGenerator U55 (G[55], P[55], X[55], Y[55]);
  GPGenerator U56 (G[56], P[56], X[56], Y[56]);
  GPGenerator U57 (G[57], P[57], X[57], Y[57]);
  GPGenerator U58 (G[58], P[58], X[58], Y[58]);
  GPGenerator U59 (G[59], P[59], X[59], Y[59]);
  GPGenerator U60 (G[60], P[60], X[60], Y[60]);
  GPGenerator U61 (G[61], P[61], X[61], Y[61]);
  GPGenerator U62 (G[62], P[62], X[62], Y[62]);
  GPGenerator U63 (G[63], P[63], X[63], Y[63]);
  CLAUnit_64 U64 (C, G, P, Cin);
endmodule

module UBZero_0_0(O);
  output [0:0] O;
  assign O[0] = 0;
endmodule

module UBCLA_15_0_63_0 (S, X, Y);
  output [64:0] S;
  input [15:0] X;
  input [63:0] Y;
  wire [63:0] Z;
  UBExtender_15_0_6000 U0 (Z[63:0], X[15:0]);
  UBPureCLA_63_0 U1 (S[64:0], Z[63:0], Y[63:0]);
endmodule

module UBCON_15_0 (O, I);
  output [15:0] O;
  input [15:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
  UB1DCON_13 U13 (O[13], I[13]);
  UB1DCON_14 U14 (O[14], I[14]);
  UB1DCON_15 U15 (O[15], I[15]);
endmodule

module UBExtender_15_0_6000 (O, I);
  output [63:0] O;
  input [15:0] I;
  UBCON_15_0 U0 (O[15:0], I[15:0]);
  UBZero_63_16 U1 (O[63:16]);
endmodule

module UBPureCLA_63_0 (S, X, Y);
  output [64:0] S;
  input [63:0] X;
  input [63:0] Y;
  wire C;
  UBPriCLA_63_0 U0 (S, X, Y, C);
  UBZero_0_0 U1 (C);
endmodule

