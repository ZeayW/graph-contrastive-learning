library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_0_0 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_0_0;

architecture UB1BPPG_0_0 of UB1BPPG_0_0 is
begin
   O <= IN1 and IN2;
end UB1BPPG_0_0;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_1_0 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_1_0;

architecture UB1BPPG_1_0 of UB1BPPG_1_0 is
begin
   O <= IN1 and IN2;
end UB1BPPG_1_0;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_2_0 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_2_0;

architecture UB1BPPG_2_0 of UB1BPPG_2_0 is
begin
   O <= IN1 and IN2;
end UB1BPPG_2_0;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_3_0 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_3_0;

architecture UB1BPPG_3_0 of UB1BPPG_3_0 is
begin
   O <= IN1 and IN2;
end UB1BPPG_3_0;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_4_0 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_4_0;

architecture UB1BPPG_4_0 of UB1BPPG_4_0 is
begin
   O <= IN1 and IN2;
end UB1BPPG_4_0;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_5_0 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_5_0;

architecture UB1BPPG_5_0 of UB1BPPG_5_0 is
begin
   O <= IN1 and IN2;
end UB1BPPG_5_0;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_6_0 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_6_0;

architecture UB1BPPG_6_0 of UB1BPPG_6_0 is
begin
   O <= IN1 and IN2;
end UB1BPPG_6_0;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_7_0 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_7_0;

architecture UB1BPPG_7_0 of UB1BPPG_7_0 is
begin
   O <= IN1 and IN2;
end UB1BPPG_7_0;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_0_1 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_0_1;

architecture UB1BPPG_0_1 of UB1BPPG_0_1 is
begin
   O <= IN1 and IN2;
end UB1BPPG_0_1;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_1_1 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_1_1;

architecture UB1BPPG_1_1 of UB1BPPG_1_1 is
begin
   O <= IN1 and IN2;
end UB1BPPG_1_1;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_2_1 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_2_1;

architecture UB1BPPG_2_1 of UB1BPPG_2_1 is
begin
   O <= IN1 and IN2;
end UB1BPPG_2_1;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_3_1 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_3_1;

architecture UB1BPPG_3_1 of UB1BPPG_3_1 is
begin
   O <= IN1 and IN2;
end UB1BPPG_3_1;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_4_1 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_4_1;

architecture UB1BPPG_4_1 of UB1BPPG_4_1 is
begin
   O <= IN1 and IN2;
end UB1BPPG_4_1;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_5_1 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_5_1;

architecture UB1BPPG_5_1 of UB1BPPG_5_1 is
begin
   O <= IN1 and IN2;
end UB1BPPG_5_1;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_6_1 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_6_1;

architecture UB1BPPG_6_1 of UB1BPPG_6_1 is
begin
   O <= IN1 and IN2;
end UB1BPPG_6_1;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_7_1 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_7_1;

architecture UB1BPPG_7_1 of UB1BPPG_7_1 is
begin
   O <= IN1 and IN2;
end UB1BPPG_7_1;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_0_2 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_0_2;

architecture UB1BPPG_0_2 of UB1BPPG_0_2 is
begin
   O <= IN1 and IN2;
end UB1BPPG_0_2;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_1_2 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_1_2;

architecture UB1BPPG_1_2 of UB1BPPG_1_2 is
begin
   O <= IN1 and IN2;
end UB1BPPG_1_2;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_2_2 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_2_2;

architecture UB1BPPG_2_2 of UB1BPPG_2_2 is
begin
   O <= IN1 and IN2;
end UB1BPPG_2_2;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_3_2 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_3_2;

architecture UB1BPPG_3_2 of UB1BPPG_3_2 is
begin
   O <= IN1 and IN2;
end UB1BPPG_3_2;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_4_2 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_4_2;

architecture UB1BPPG_4_2 of UB1BPPG_4_2 is
begin
   O <= IN1 and IN2;
end UB1BPPG_4_2;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_5_2 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_5_2;

architecture UB1BPPG_5_2 of UB1BPPG_5_2 is
begin
   O <= IN1 and IN2;
end UB1BPPG_5_2;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_6_2 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_6_2;

architecture UB1BPPG_6_2 of UB1BPPG_6_2 is
begin
   O <= IN1 and IN2;
end UB1BPPG_6_2;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_7_2 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_7_2;

architecture UB1BPPG_7_2 of UB1BPPG_7_2 is
begin
   O <= IN1 and IN2;
end UB1BPPG_7_2;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_0_3 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_0_3;

architecture UB1BPPG_0_3 of UB1BPPG_0_3 is
begin
   O <= IN1 and IN2;
end UB1BPPG_0_3;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_1_3 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_1_3;

architecture UB1BPPG_1_3 of UB1BPPG_1_3 is
begin
   O <= IN1 and IN2;
end UB1BPPG_1_3;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_2_3 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_2_3;

architecture UB1BPPG_2_3 of UB1BPPG_2_3 is
begin
   O <= IN1 and IN2;
end UB1BPPG_2_3;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_3_3 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_3_3;

architecture UB1BPPG_3_3 of UB1BPPG_3_3 is
begin
   O <= IN1 and IN2;
end UB1BPPG_3_3;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_4_3 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_4_3;

architecture UB1BPPG_4_3 of UB1BPPG_4_3 is
begin
   O <= IN1 and IN2;
end UB1BPPG_4_3;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_5_3 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_5_3;

architecture UB1BPPG_5_3 of UB1BPPG_5_3 is
begin
   O <= IN1 and IN2;
end UB1BPPG_5_3;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_6_3 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_6_3;

architecture UB1BPPG_6_3 of UB1BPPG_6_3 is
begin
   O <= IN1 and IN2;
end UB1BPPG_6_3;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_7_3 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_7_3;

architecture UB1BPPG_7_3 of UB1BPPG_7_3 is
begin
   O <= IN1 and IN2;
end UB1BPPG_7_3;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_0_4 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_0_4;

architecture UB1BPPG_0_4 of UB1BPPG_0_4 is
begin
   O <= IN1 and IN2;
end UB1BPPG_0_4;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_1_4 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_1_4;

architecture UB1BPPG_1_4 of UB1BPPG_1_4 is
begin
   O <= IN1 and IN2;
end UB1BPPG_1_4;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_2_4 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_2_4;

architecture UB1BPPG_2_4 of UB1BPPG_2_4 is
begin
   O <= IN1 and IN2;
end UB1BPPG_2_4;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_3_4 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_3_4;

architecture UB1BPPG_3_4 of UB1BPPG_3_4 is
begin
   O <= IN1 and IN2;
end UB1BPPG_3_4;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_4_4 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_4_4;

architecture UB1BPPG_4_4 of UB1BPPG_4_4 is
begin
   O <= IN1 and IN2;
end UB1BPPG_4_4;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_5_4 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_5_4;

architecture UB1BPPG_5_4 of UB1BPPG_5_4 is
begin
   O <= IN1 and IN2;
end UB1BPPG_5_4;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_6_4 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_6_4;

architecture UB1BPPG_6_4 of UB1BPPG_6_4 is
begin
   O <= IN1 and IN2;
end UB1BPPG_6_4;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_7_4 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_7_4;

architecture UB1BPPG_7_4 of UB1BPPG_7_4 is
begin
   O <= IN1 and IN2;
end UB1BPPG_7_4;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_0_5 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_0_5;

architecture UB1BPPG_0_5 of UB1BPPG_0_5 is
begin
   O <= IN1 and IN2;
end UB1BPPG_0_5;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_1_5 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_1_5;

architecture UB1BPPG_1_5 of UB1BPPG_1_5 is
begin
   O <= IN1 and IN2;
end UB1BPPG_1_5;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_2_5 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_2_5;

architecture UB1BPPG_2_5 of UB1BPPG_2_5 is
begin
   O <= IN1 and IN2;
end UB1BPPG_2_5;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_3_5 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_3_5;

architecture UB1BPPG_3_5 of UB1BPPG_3_5 is
begin
   O <= IN1 and IN2;
end UB1BPPG_3_5;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_4_5 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_4_5;

architecture UB1BPPG_4_5 of UB1BPPG_4_5 is
begin
   O <= IN1 and IN2;
end UB1BPPG_4_5;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_5_5 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_5_5;

architecture UB1BPPG_5_5 of UB1BPPG_5_5 is
begin
   O <= IN1 and IN2;
end UB1BPPG_5_5;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_6_5 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_6_5;

architecture UB1BPPG_6_5 of UB1BPPG_6_5 is
begin
   O <= IN1 and IN2;
end UB1BPPG_6_5;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_7_5 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_7_5;

architecture UB1BPPG_7_5 of UB1BPPG_7_5 is
begin
   O <= IN1 and IN2;
end UB1BPPG_7_5;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_0_6 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_0_6;

architecture UB1BPPG_0_6 of UB1BPPG_0_6 is
begin
   O <= IN1 and IN2;
end UB1BPPG_0_6;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_1_6 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_1_6;

architecture UB1BPPG_1_6 of UB1BPPG_1_6 is
begin
   O <= IN1 and IN2;
end UB1BPPG_1_6;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_2_6 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_2_6;

architecture UB1BPPG_2_6 of UB1BPPG_2_6 is
begin
   O <= IN1 and IN2;
end UB1BPPG_2_6;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_3_6 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_3_6;

architecture UB1BPPG_3_6 of UB1BPPG_3_6 is
begin
   O <= IN1 and IN2;
end UB1BPPG_3_6;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_4_6 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_4_6;

architecture UB1BPPG_4_6 of UB1BPPG_4_6 is
begin
   O <= IN1 and IN2;
end UB1BPPG_4_6;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_5_6 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_5_6;

architecture UB1BPPG_5_6 of UB1BPPG_5_6 is
begin
   O <= IN1 and IN2;
end UB1BPPG_5_6;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_6_6 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_6_6;

architecture UB1BPPG_6_6 of UB1BPPG_6_6 is
begin
   O <= IN1 and IN2;
end UB1BPPG_6_6;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_7_6 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_7_6;

architecture UB1BPPG_7_6 of UB1BPPG_7_6 is
begin
   O <= IN1 and IN2;
end UB1BPPG_7_6;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_0_7 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_0_7;

architecture UB1BPPG_0_7 of UB1BPPG_0_7 is
begin
   O <= IN1 and IN2;
end UB1BPPG_0_7;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_1_7 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_1_7;

architecture UB1BPPG_1_7 of UB1BPPG_1_7 is
begin
   O <= IN1 and IN2;
end UB1BPPG_1_7;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_2_7 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_2_7;

architecture UB1BPPG_2_7 of UB1BPPG_2_7 is
begin
   O <= IN1 and IN2;
end UB1BPPG_2_7;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_3_7 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_3_7;

architecture UB1BPPG_3_7 of UB1BPPG_3_7 is
begin
   O <= IN1 and IN2;
end UB1BPPG_3_7;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_4_7 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_4_7;

architecture UB1BPPG_4_7 of UB1BPPG_4_7 is
begin
   O <= IN1 and IN2;
end UB1BPPG_4_7;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_5_7 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_5_7;

architecture UB1BPPG_5_7 of UB1BPPG_5_7 is
begin
   O <= IN1 and IN2;
end UB1BPPG_5_7;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_6_7 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_6_7;

architecture UB1BPPG_6_7 of UB1BPPG_6_7 is
begin
   O <= IN1 and IN2;
end UB1BPPG_6_7;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1BPPG_7_7 is
  port ( O : out std_logic;
         IN1 : in  std_logic;
         IN2 : in  std_logic );
end UB1BPPG_7_7;

architecture UB1BPPG_7_7 of UB1BPPG_7_7 is
begin
   O <= IN1 and IN2;
end UB1BPPG_7_7;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1DCON_0 is
  port ( O : out std_logic;
         I : in  std_logic );
end UB1DCON_0;

architecture UB1DCON_0 of UB1DCON_0 is
begin
   O <= I;
end UB1DCON_0;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBHA_1 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic );
end UBHA_1;

architecture UBHA_1 of UBHA_1 is
begin
   C <= X and Y;
   S <= X xor Y;
end UBHA_1;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBFA_2 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic;
         Z : in  std_logic );
end UBFA_2;

architecture UBFA_2 of UBFA_2 is
begin
   C <= ( X and Y ) or ( Y and Z ) or ( Z and X );
   S <= X xor Y xor Z;
end UBFA_2;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBFA_3 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic;
         Z : in  std_logic );
end UBFA_3;

architecture UBFA_3 of UBFA_3 is
begin
   C <= ( X and Y ) or ( Y and Z ) or ( Z and X );
   S <= X xor Y xor Z;
end UBFA_3;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBFA_4 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic;
         Z : in  std_logic );
end UBFA_4;

architecture UBFA_4 of UBFA_4 is
begin
   C <= ( X and Y ) or ( Y and Z ) or ( Z and X );
   S <= X xor Y xor Z;
end UBFA_4;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBFA_5 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic;
         Z : in  std_logic );
end UBFA_5;

architecture UBFA_5 of UBFA_5 is
begin
   C <= ( X and Y ) or ( Y and Z ) or ( Z and X );
   S <= X xor Y xor Z;
end UBFA_5;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBFA_6 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic;
         Z : in  std_logic );
end UBFA_6;

architecture UBFA_6 of UBFA_6 is
begin
   C <= ( X and Y ) or ( Y and Z ) or ( Z and X );
   S <= X xor Y xor Z;
end UBFA_6;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBFA_7 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic;
         Z : in  std_logic );
end UBFA_7;

architecture UBFA_7 of UBFA_7 is
begin
   C <= ( X and Y ) or ( Y and Z ) or ( Z and X );
   S <= X xor Y xor Z;
end UBFA_7;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBHA_8 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic );
end UBHA_8;

architecture UBHA_8 of UBHA_8 is
begin
   C <= X and Y;
   S <= X xor Y;
end UBHA_8;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1DCON_9 is
  port ( O : out std_logic;
         I : in  std_logic );
end UB1DCON_9;

architecture UB1DCON_9 of UB1DCON_9 is
begin
   O <= I;
end UB1DCON_9;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1DCON_1 is
  port ( O : out std_logic;
         I : in  std_logic );
end UB1DCON_1;

architecture UB1DCON_1 of UB1DCON_1 is
begin
   O <= I;
end UB1DCON_1;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBHA_2 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic );
end UBHA_2;

architecture UBHA_2 of UBHA_2 is
begin
   C <= X and Y;
   S <= X xor Y;
end UBHA_2;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBFA_8 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic;
         Z : in  std_logic );
end UBFA_8;

architecture UBFA_8 of UBFA_8 is
begin
   C <= ( X and Y ) or ( Y and Z ) or ( Z and X );
   S <= X xor Y xor Z;
end UBFA_8;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBFA_9 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic;
         Z : in  std_logic );
end UBFA_9;

architecture UBFA_9 of UBFA_9 is
begin
   C <= ( X and Y ) or ( Y and Z ) or ( Z and X );
   S <= X xor Y xor Z;
end UBFA_9;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1DCON_10 is
  port ( O : out std_logic;
         I : in  std_logic );
end UB1DCON_10;

architecture UB1DCON_10 of UB1DCON_10 is
begin
   O <= I;
end UB1DCON_10;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1DCON_2 is
  port ( O : out std_logic;
         I : in  std_logic );
end UB1DCON_2;

architecture UB1DCON_2 of UB1DCON_2 is
begin
   O <= I;
end UB1DCON_2;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBHA_3 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic );
end UBHA_3;

architecture UBHA_3 of UBHA_3 is
begin
   C <= X and Y;
   S <= X xor Y;
end UBHA_3;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBFA_10 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic;
         Z : in  std_logic );
end UBFA_10;

architecture UBFA_10 of UBFA_10 is
begin
   C <= ( X and Y ) or ( Y and Z ) or ( Z and X );
   S <= X xor Y xor Z;
end UBFA_10;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1DCON_11 is
  port ( O : out std_logic;
         I : in  std_logic );
end UB1DCON_11;

architecture UB1DCON_11 of UB1DCON_11 is
begin
   O <= I;
end UB1DCON_11;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1DCON_3 is
  port ( O : out std_logic;
         I : in  std_logic );
end UB1DCON_3;

architecture UB1DCON_3 of UB1DCON_3 is
begin
   O <= I;
end UB1DCON_3;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBHA_4 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic );
end UBHA_4;

architecture UBHA_4 of UBHA_4 is
begin
   C <= X and Y;
   S <= X xor Y;
end UBHA_4;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBFA_11 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic;
         Z : in  std_logic );
end UBFA_11;

architecture UBFA_11 of UBFA_11 is
begin
   C <= ( X and Y ) or ( Y and Z ) or ( Z and X );
   S <= X xor Y xor Z;
end UBFA_11;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1DCON_12 is
  port ( O : out std_logic;
         I : in  std_logic );
end UB1DCON_12;

architecture UB1DCON_12 of UB1DCON_12 is
begin
   O <= I;
end UB1DCON_12;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1DCON_4 is
  port ( O : out std_logic;
         I : in  std_logic );
end UB1DCON_4;

architecture UB1DCON_4 of UB1DCON_4 is
begin
   O <= I;
end UB1DCON_4;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBHA_5 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic );
end UBHA_5;

architecture UBHA_5 of UBHA_5 is
begin
   C <= X and Y;
   S <= X xor Y;
end UBHA_5;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBFA_12 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic;
         Z : in  std_logic );
end UBFA_12;

architecture UBFA_12 of UBFA_12 is
begin
   C <= ( X and Y ) or ( Y and Z ) or ( Z and X );
   S <= X xor Y xor Z;
end UBFA_12;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1DCON_13 is
  port ( O : out std_logic;
         I : in  std_logic );
end UB1DCON_13;

architecture UB1DCON_13 of UB1DCON_13 is
begin
   O <= I;
end UB1DCON_13;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1DCON_5 is
  port ( O : out std_logic;
         I : in  std_logic );
end UB1DCON_5;

architecture UB1DCON_5 of UB1DCON_5 is
begin
   O <= I;
end UB1DCON_5;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBHA_6 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic );
end UBHA_6;

architecture UBHA_6 of UBHA_6 is
begin
   C <= X and Y;
   S <= X xor Y;
end UBHA_6;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBFA_13 is
  port ( C : out std_logic;
         S : out std_logic;
         X : in  std_logic;
         Y : in  std_logic;
         Z : in  std_logic );
end UBFA_13;

architecture UBFA_13 of UBFA_13 is
begin
   C <= ( X and Y ) or ( Y and Z ) or ( Z and X );
   S <= X xor Y xor Z;
end UBFA_13;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1DCON_14 is
  port ( O : out std_logic;
         I : in  std_logic );
end UB1DCON_14;

architecture UB1DCON_14 of UB1DCON_14 is
begin
   O <= I;
end UB1DCON_14;

library IEEE;
use IEEE.std_logic_1164.all;

entity GPGenerator is
  port ( Go : out std_logic;
         Po : out std_logic;
         A : in  std_logic;
         B : in  std_logic );
end GPGenerator;

architecture GPGenerator of GPGenerator is
begin
   Go <= A and B;
   Po <= A xor B;
end GPGenerator;

library IEEE;
use IEEE.std_logic_1164.all;

entity CLAUnit_8 is
  port ( C : out std_logic_vector ( 8 downto 1 );
         G : in  std_logic_vector ( 7 downto 0 );
         P : in  std_logic_vector ( 7 downto 0 );
         Cin : in  std_logic );
end CLAUnit_8;

architecture CLAUnit_8 of CLAUnit_8 is
begin
   C(1) <= G(0) or ( P(0) and Cin );
   C(2) <= G(1) or ( P(1) and G(0) ) or ( P(1) and P(0) and Cin );
   C(3) <= G(2) or ( P(2) and G(1) ) or ( P(2) and P(1) and G(0) ) or ( P(2) and P(1) and P(0) and Cin );
   C(4) <= G(3) or ( P(3) and G(2) ) or ( P(3) and P(2) and G(1) ) or ( P(3) and P(2) and P(1) and G(0) ) or ( P(3) and P(2) and P(1) and P(0) and Cin );
   C(5) <= G(4) or ( P(4) and G(3) ) or ( P(4) and P(3) and G(2) ) or ( P(4) and P(3) and P(2) and G(1) ) or ( P(4) and P(3) and P(2) and P(1) and G(0) ) or ( P(4) and P(3) and P(2) and P(1) and P(0) and
 Cin );
   C(6) <= G(5) or ( P(5) and G(4) ) or ( P(5) and P(4) and G(3) ) or ( P(5) and P(4) and P(3) and G(2) ) or ( P(5) and P(4) and P(3) and P(2) and G(1) ) or ( P(5) and P(4) and P(3) and P(2) and P(1) and
 G(0) ) or ( P(5) and P(4) and P(3) and P(2) and P(1) and P(0) and Cin );
   C(7) <= G(6) or ( P(6) and G(5) ) or ( P(6) and P(5) and G(4) ) or ( P(6) and P(5) and P(4) and G(3) ) or ( P(6) and P(5) and P(4) and P(3) and G(2) ) or ( P(6) and P(5) and P(4) and P(3) and P(2) and
 G(1) ) or ( P(6) and P(5) and P(4) and P(3) and P(2) and P(1) and G(0) ) or ( P(6) and P(5) and P(4) and P(3) and P(2) and P(1) and P(0) and Cin );
   C(8) <= G(7) or ( P(7) and G(6) ) or ( P(7) and P(6) and G(5) ) or ( P(7) and P(6) and P(5) and G(4) ) or ( P(7) and P(6) and P(5) and P(4) and G(3) ) or ( P(7) and P(6) and P(5) and P(4) and P(3) and
 G(2) ) or ( P(7) and P(6) and P(5) and P(4) and P(3) and P(2) and G(1) ) or ( P(7) and P(6) and P(5) and P(4) and P(3) and P(2) and P(1) and G(0) ) or ( P(7) and P(6) and P(5) and P(4) and P(3) and P(2)
 and P(1) and P(0) and Cin );
end CLAUnit_8;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBPriCLA_14_7 is
  port ( S : out std_logic_vector ( 15 downto 7 );
         X : in  std_logic_vector ( 14 downto 7 );
         Y : in  std_logic_vector ( 14 downto 7 );
         Cin : in  std_logic );
end UBPriCLA_14_7;

architecture UBPriCLA_14_7 of UBPriCLA_14_7 is
  component GPGenerator
    port ( Go : out std_logic;
           Po : out std_logic;
           A : in  std_logic;
           B : in  std_logic );
  end component;
  component CLAUnit_8
    port ( C : out std_logic_vector ( 8 downto 1 );
           G : in  std_logic_vector ( 7 downto 0 );
           P : in  std_logic_vector ( 7 downto 0 );
           Cin : in  std_logic );
  end component;
  signal C :  std_logic_vector ( 15 downto 8 );
  signal G :  std_logic_vector ( 14 downto 7 );
  signal P :  std_logic_vector ( 14 downto 7 );
begin
   S(7) <= Cin xor P(7);
   S(8) <= C(8) xor P(8);
   S(9) <= C(9) xor P(9);
   S(10) <= C(10) xor P(10);
   S(11) <= C(11) xor P(11);
   S(12) <= C(12) xor P(12);
   S(13) <= C(13) xor P(13);
   S(14) <= C(14) xor P(14);
   S(15) <= C(15);
  U0:GPGenerator port map (G(7), P(7), X(7), Y(7));
  U1:GPGenerator port map (G(8), P(8), X(8), Y(8));
  U2:GPGenerator port map (G(9), P(9), X(9), Y(9));
  U3:GPGenerator port map (G(10), P(10), X(10)
, Y(10));
  U4:GPGenerator port map (G(11), P(11), X(11), Y(11));
  U5:GPGenerator port map (G(12), P(12), X(12), Y(12));
  U6:GPGenerator port map (G(13), P(13), X(13), Y(13));
  U7:GPGenerator port map (
G(14), P(14), X(14), Y(14));
  U8:CLAUnit_8 port map (C, G, P, Cin);
end UBPriCLA_14_7;

library IEEE;
use IEEE.std_logic_1164.all;

entity UBZero_7_7 is
  port ( O : out std_logic );
end UBZero_7_7;

architecture UBZero_7_7 of UBZero_7_7 is
begin
   O <= '0';
end UBZero_7_7;

library IEEE;
use IEEE.std_logic_1164.all;

entity UB1DCON_6 is
  port ( O : out std_logic;
         I : in  std_logic );
end UB1DCON_6;

architecture UB1DCON_6 of UB1DCON_6 is
begin
   O <= I;
end UB1DCON_6;

library IEEE;
use IEEE.std_logic_1164.all;

entity Multiplier_7_0_7_000 is
  port ( P : out std_logic_vector ( 15 downto 0 );
         IN1 : in  std_logic_vector ( 7 downto 0 );
         IN2 : in  std_logic_vector ( 7 downto 0 ) );
end Multiplier_7_0_7_000;

architecture Multiplier_7_0_7_000 of Multiplier_7_0_7_000 is
  component MultUB_STD_ARY_CL000
    port ( P : out std_logic_vector ( 15 downto 0 );
           IN1 : in  std_logic_vector ( 7 downto 0 );
           IN2 : in  std_logic_vector ( 7 downto 0 ) );
  end component;
  signal W :  std_logic_vector ( 15 downto 0 );
begin
   P(0) <= W(0);
   P(1) <= W(1);
   P(2) <= W(2);
   P(3) <= W(3);
   P(4) <= W(4);
   P(5) <= W(5);
   P(6) <= W(6);
   P(7) <= W(7);
   P(8) <= W(8);
   P(9) <= W(9);
   P(10) <= W(10);
   P(11) <= W(11);
   P(12) <= W(12);
   P(13) <= W(13);
   P(14) <= W(14);
   P(15) <= W(15);
  U0:MultUB_STD_ARY_CL000 port map (W, IN1, IN2);
end Multiplier_7_0_7_000;

