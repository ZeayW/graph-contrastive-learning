/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: UBKSA_31_0_47_0

  Operand-1 length: 32
  Operand-2 length: 48
  Two-operand addition algorithm: Kogge-Stone adder
----------------------------------------------------------------------------*/

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_21(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_23(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_24(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_25(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_27(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_28(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_29(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_30(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_31(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_47_32(O);
  output [47:32] O;
  assign O[32] = 0;
  assign O[33] = 0;
  assign O[34] = 0;
  assign O[35] = 0;
  assign O[36] = 0;
  assign O[37] = 0;
  assign O[38] = 0;
  assign O[39] = 0;
  assign O[40] = 0;
  assign O[41] = 0;
  assign O[42] = 0;
  assign O[43] = 0;
  assign O[44] = 0;
  assign O[45] = 0;
  assign O[46] = 0;
  assign O[47] = 0;
endmodule

module GPGenerator(Go, Po, A, B);
  output Go;
  output Po;
  input A;
  input B;
  assign Go = A & B;
  assign Po = A ^ B;
endmodule

module CarryOperator(Go, Po, Gi1, Pi1, Gi2, Pi2);
  output Go;
  output Po;
  input Gi1;
  input Gi2;
  input Pi1;
  input Pi2;
  assign Go = Gi1 | ( Gi2 & Pi1 );
  assign Po = Pi1 & Pi2;
endmodule

module UBPriKSA_47_0(S, X, Y, Cin);
  output [48:0] S;
  input Cin;
  input [47:0] X;
  input [47:0] Y;
  wire [47:0] G0;
  wire [47:0] G1;
  wire [47:0] G2;
  wire [47:0] G3;
  wire [47:0] G4;
  wire [47:0] G5;
  wire [47:0] G6;
  wire [47:0] P0;
  wire [47:0] P1;
  wire [47:0] P2;
  wire [47:0] P3;
  wire [47:0] P4;
  wire [47:0] P5;
  wire [47:0] P6;
  assign P1[0] = P0[0];
  assign G1[0] = G0[0];
  assign P2[0] = P1[0];
  assign G2[0] = G1[0];
  assign P2[1] = P1[1];
  assign G2[1] = G1[1];
  assign P3[0] = P2[0];
  assign G3[0] = G2[0];
  assign P3[1] = P2[1];
  assign G3[1] = G2[1];
  assign P3[2] = P2[2];
  assign G3[2] = G2[2];
  assign P3[3] = P2[3];
  assign G3[3] = G2[3];
  assign P4[0] = P3[0];
  assign G4[0] = G3[0];
  assign P4[1] = P3[1];
  assign G4[1] = G3[1];
  assign P4[2] = P3[2];
  assign G4[2] = G3[2];
  assign P4[3] = P3[3];
  assign G4[3] = G3[3];
  assign P4[4] = P3[4];
  assign G4[4] = G3[4];
  assign P4[5] = P3[5];
  assign G4[5] = G3[5];
  assign P4[6] = P3[6];
  assign G4[6] = G3[6];
  assign P4[7] = P3[7];
  assign G4[7] = G3[7];
  assign P5[0] = P4[0];
  assign G5[0] = G4[0];
  assign P5[1] = P4[1];
  assign G5[1] = G4[1];
  assign P5[2] = P4[2];
  assign G5[2] = G4[2];
  assign P5[3] = P4[3];
  assign G5[3] = G4[3];
  assign P5[4] = P4[4];
  assign G5[4] = G4[4];
  assign P5[5] = P4[5];
  assign G5[5] = G4[5];
  assign P5[6] = P4[6];
  assign G5[6] = G4[6];
  assign P5[7] = P4[7];
  assign G5[7] = G4[7];
  assign P5[8] = P4[8];
  assign G5[8] = G4[8];
  assign P5[9] = P4[9];
  assign G5[9] = G4[9];
  assign P5[10] = P4[10];
  assign G5[10] = G4[10];
  assign P5[11] = P4[11];
  assign G5[11] = G4[11];
  assign P5[12] = P4[12];
  assign G5[12] = G4[12];
  assign P5[13] = P4[13];
  assign G5[13] = G4[13];
  assign P5[14] = P4[14];
  assign G5[14] = G4[14];
  assign P5[15] = P4[15];
  assign G5[15] = G4[15];
  assign P6[0] = P5[0];
  assign G6[0] = G5[0];
  assign P6[1] = P5[1];
  assign G6[1] = G5[1];
  assign P6[2] = P5[2];
  assign G6[2] = G5[2];
  assign P6[3] = P5[3];
  assign G6[3] = G5[3];
  assign P6[4] = P5[4];
  assign G6[4] = G5[4];
  assign P6[5] = P5[5];
  assign G6[5] = G5[5];
  assign P6[6] = P5[6];
  assign G6[6] = G5[6];
  assign P6[7] = P5[7];
  assign G6[7] = G5[7];
  assign P6[8] = P5[8];
  assign G6[8] = G5[8];
  assign P6[9] = P5[9];
  assign G6[9] = G5[9];
  assign P6[10] = P5[10];
  assign G6[10] = G5[10];
  assign P6[11] = P5[11];
  assign G6[11] = G5[11];
  assign P6[12] = P5[12];
  assign G6[12] = G5[12];
  assign P6[13] = P5[13];
  assign G6[13] = G5[13];
  assign P6[14] = P5[14];
  assign G6[14] = G5[14];
  assign P6[15] = P5[15];
  assign G6[15] = G5[15];
  assign P6[16] = P5[16];
  assign G6[16] = G5[16];
  assign P6[17] = P5[17];
  assign G6[17] = G5[17];
  assign P6[18] = P5[18];
  assign G6[18] = G5[18];
  assign P6[19] = P5[19];
  assign G6[19] = G5[19];
  assign P6[20] = P5[20];
  assign G6[20] = G5[20];
  assign P6[21] = P5[21];
  assign G6[21] = G5[21];
  assign P6[22] = P5[22];
  assign G6[22] = G5[22];
  assign P6[23] = P5[23];
  assign G6[23] = G5[23];
  assign P6[24] = P5[24];
  assign G6[24] = G5[24];
  assign P6[25] = P5[25];
  assign G6[25] = G5[25];
  assign P6[26] = P5[26];
  assign G6[26] = G5[26];
  assign P6[27] = P5[27];
  assign G6[27] = G5[27];
  assign P6[28] = P5[28];
  assign G6[28] = G5[28];
  assign P6[29] = P5[29];
  assign G6[29] = G5[29];
  assign P6[30] = P5[30];
  assign G6[30] = G5[30];
  assign P6[31] = P5[31];
  assign G6[31] = G5[31];
  assign S[0] = Cin ^ P0[0];
  assign S[1] = ( G6[0] | ( P6[0] & Cin ) ) ^ P0[1];
  assign S[2] = ( G6[1] | ( P6[1] & Cin ) ) ^ P0[2];
  assign S[3] = ( G6[2] | ( P6[2] & Cin ) ) ^ P0[3];
  assign S[4] = ( G6[3] | ( P6[3] & Cin ) ) ^ P0[4];
  assign S[5] = ( G6[4] | ( P6[4] & Cin ) ) ^ P0[5];
  assign S[6] = ( G6[5] | ( P6[5] & Cin ) ) ^ P0[6];
  assign S[7] = ( G6[6] | ( P6[6] & Cin ) ) ^ P0[7];
  assign S[8] = ( G6[7] | ( P6[7] & Cin ) ) ^ P0[8];
  assign S[9] = ( G6[8] | ( P6[8] & Cin ) ) ^ P0[9];
  assign S[10] = ( G6[9] | ( P6[9] & Cin ) ) ^ P0[10];
  assign S[11] = ( G6[10] | ( P6[10] & Cin ) ) ^ P0[11];
  assign S[12] = ( G6[11] | ( P6[11] & Cin ) ) ^ P0[12];
  assign S[13] = ( G6[12] | ( P6[12] & Cin ) ) ^ P0[13];
  assign S[14] = ( G6[13] | ( P6[13] & Cin ) ) ^ P0[14];
  assign S[15] = ( G6[14] | ( P6[14] & Cin ) ) ^ P0[15];
  assign S[16] = ( G6[15] | ( P6[15] & Cin ) ) ^ P0[16];
  assign S[17] = ( G6[16] | ( P6[16] & Cin ) ) ^ P0[17];
  assign S[18] = ( G6[17] | ( P6[17] & Cin ) ) ^ P0[18];
  assign S[19] = ( G6[18] | ( P6[18] & Cin ) ) ^ P0[19];
  assign S[20] = ( G6[19] | ( P6[19] & Cin ) ) ^ P0[20];
  assign S[21] = ( G6[20] | ( P6[20] & Cin ) ) ^ P0[21];
  assign S[22] = ( G6[21] | ( P6[21] & Cin ) ) ^ P0[22];
  assign S[23] = ( G6[22] | ( P6[22] & Cin ) ) ^ P0[23];
  assign S[24] = ( G6[23] | ( P6[23] & Cin ) ) ^ P0[24];
  assign S[25] = ( G6[24] | ( P6[24] & Cin ) ) ^ P0[25];
  assign S[26] = ( G6[25] | ( P6[25] & Cin ) ) ^ P0[26];
  assign S[27] = ( G6[26] | ( P6[26] & Cin ) ) ^ P0[27];
  assign S[28] = ( G6[27] | ( P6[27] & Cin ) ) ^ P0[28];
  assign S[29] = ( G6[28] | ( P6[28] & Cin ) ) ^ P0[29];
  assign S[30] = ( G6[29] | ( P6[29] & Cin ) ) ^ P0[30];
  assign S[31] = ( G6[30] | ( P6[30] & Cin ) ) ^ P0[31];
  assign S[32] = ( G6[31] | ( P6[31] & Cin ) ) ^ P0[32];
  assign S[33] = ( G6[32] | ( P6[32] & Cin ) ) ^ P0[33];
  assign S[34] = ( G6[33] | ( P6[33] & Cin ) ) ^ P0[34];
  assign S[35] = ( G6[34] | ( P6[34] & Cin ) ) ^ P0[35];
  assign S[36] = ( G6[35] | ( P6[35] & Cin ) ) ^ P0[36];
  assign S[37] = ( G6[36] | ( P6[36] & Cin ) ) ^ P0[37];
  assign S[38] = ( G6[37] | ( P6[37] & Cin ) ) ^ P0[38];
  assign S[39] = ( G6[38] | ( P6[38] & Cin ) ) ^ P0[39];
  assign S[40] = ( G6[39] | ( P6[39] & Cin ) ) ^ P0[40];
  assign S[41] = ( G6[40] | ( P6[40] & Cin ) ) ^ P0[41];
  assign S[42] = ( G6[41] | ( P6[41] & Cin ) ) ^ P0[42];
  assign S[43] = ( G6[42] | ( P6[42] & Cin ) ) ^ P0[43];
  assign S[44] = ( G6[43] | ( P6[43] & Cin ) ) ^ P0[44];
  assign S[45] = ( G6[44] | ( P6[44] & Cin ) ) ^ P0[45];
  assign S[46] = ( G6[45] | ( P6[45] & Cin ) ) ^ P0[46];
  assign S[47] = ( G6[46] | ( P6[46] & Cin ) ) ^ P0[47];
  assign S[48] = G6[47] | ( P6[47] & Cin );
  GPGenerator U0 (G0[0], P0[0], X[0], Y[0]);
  GPGenerator U1 (G0[1], P0[1], X[1], Y[1]);
  GPGenerator U2 (G0[2], P0[2], X[2], Y[2]);
  GPGenerator U3 (G0[3], P0[3], X[3], Y[3]);
  GPGenerator U4 (G0[4], P0[4], X[4], Y[4]);
  GPGenerator U5 (G0[5], P0[5], X[5], Y[5]);
  GPGenerator U6 (G0[6], P0[6], X[6], Y[6]);
  GPGenerator U7 (G0[7], P0[7], X[7], Y[7]);
  GPGenerator U8 (G0[8], P0[8], X[8], Y[8]);
  GPGenerator U9 (G0[9], P0[9], X[9], Y[9]);
  GPGenerator U10 (G0[10], P0[10], X[10], Y[10]);
  GPGenerator U11 (G0[11], P0[11], X[11], Y[11]);
  GPGenerator U12 (G0[12], P0[12], X[12], Y[12]);
  GPGenerator U13 (G0[13], P0[13], X[13], Y[13]);
  GPGenerator U14 (G0[14], P0[14], X[14], Y[14]);
  GPGenerator U15 (G0[15], P0[15], X[15], Y[15]);
  GPGenerator U16 (G0[16], P0[16], X[16], Y[16]);
  GPGenerator U17 (G0[17], P0[17], X[17], Y[17]);
  GPGenerator U18 (G0[18], P0[18], X[18], Y[18]);
  GPGenerator U19 (G0[19], P0[19], X[19], Y[19]);
  GPGenerator U20 (G0[20], P0[20], X[20], Y[20]);
  GPGenerator U21 (G0[21], P0[21], X[21], Y[21]);
  GPGenerator U22 (G0[22], P0[22], X[22], Y[22]);
  GPGenerator U23 (G0[23], P0[23], X[23], Y[23]);
  GPGenerator U24 (G0[24], P0[24], X[24], Y[24]);
  GPGenerator U25 (G0[25], P0[25], X[25], Y[25]);
  GPGenerator U26 (G0[26], P0[26], X[26], Y[26]);
  GPGenerator U27 (G0[27], P0[27], X[27], Y[27]);
  GPGenerator U28 (G0[28], P0[28], X[28], Y[28]);
  GPGenerator U29 (G0[29], P0[29], X[29], Y[29]);
  GPGenerator U30 (G0[30], P0[30], X[30], Y[30]);
  GPGenerator U31 (G0[31], P0[31], X[31], Y[31]);
  GPGenerator U32 (G0[32], P0[32], X[32], Y[32]);
  GPGenerator U33 (G0[33], P0[33], X[33], Y[33]);
  GPGenerator U34 (G0[34], P0[34], X[34], Y[34]);
  GPGenerator U35 (G0[35], P0[35], X[35], Y[35]);
  GPGenerator U36 (G0[36], P0[36], X[36], Y[36]);
  GPGenerator U37 (G0[37], P0[37], X[37], Y[37]);
  GPGenerator U38 (G0[38], P0[38], X[38], Y[38]);
  GPGenerator U39 (G0[39], P0[39], X[39], Y[39]);
  GPGenerator U40 (G0[40], P0[40], X[40], Y[40]);
  GPGenerator U41 (G0[41], P0[41], X[41], Y[41]);
  GPGenerator U42 (G0[42], P0[42], X[42], Y[42]);
  GPGenerator U43 (G0[43], P0[43], X[43], Y[43]);
  GPGenerator U44 (G0[44], P0[44], X[44], Y[44]);
  GPGenerator U45 (G0[45], P0[45], X[45], Y[45]);
  GPGenerator U46 (G0[46], P0[46], X[46], Y[46]);
  GPGenerator U47 (G0[47], P0[47], X[47], Y[47]);
  CarryOperator U48 (G1[1], P1[1], G0[1], P0[1], G0[0], P0[0]);
  CarryOperator U49 (G1[2], P1[2], G0[2], P0[2], G0[1], P0[1]);
  CarryOperator U50 (G1[3], P1[3], G0[3], P0[3], G0[2], P0[2]);
  CarryOperator U51 (G1[4], P1[4], G0[4], P0[4], G0[3], P0[3]);
  CarryOperator U52 (G1[5], P1[5], G0[5], P0[5], G0[4], P0[4]);
  CarryOperator U53 (G1[6], P1[6], G0[6], P0[6], G0[5], P0[5]);
  CarryOperator U54 (G1[7], P1[7], G0[7], P0[7], G0[6], P0[6]);
  CarryOperator U55 (G1[8], P1[8], G0[8], P0[8], G0[7], P0[7]);
  CarryOperator U56 (G1[9], P1[9], G0[9], P0[9], G0[8], P0[8]);
  CarryOperator U57 (G1[10], P1[10], G0[10], P0[10], G0[9], P0[9]);
  CarryOperator U58 (G1[11], P1[11], G0[11], P0[11], G0[10], P0[10]);
  CarryOperator U59 (G1[12], P1[12], G0[12], P0[12], G0[11], P0[11]);
  CarryOperator U60 (G1[13], P1[13], G0[13], P0[13], G0[12], P0[12]);
  CarryOperator U61 (G1[14], P1[14], G0[14], P0[14], G0[13], P0[13]);
  CarryOperator U62 (G1[15], P1[15], G0[15], P0[15], G0[14], P0[14]);
  CarryOperator U63 (G1[16], P1[16], G0[16], P0[16], G0[15], P0[15]);
  CarryOperator U64 (G1[17], P1[17], G0[17], P0[17], G0[16], P0[16]);
  CarryOperator U65 (G1[18], P1[18], G0[18], P0[18], G0[17], P0[17]);
  CarryOperator U66 (G1[19], P1[19], G0[19], P0[19], G0[18], P0[18]);
  CarryOperator U67 (G1[20], P1[20], G0[20], P0[20], G0[19], P0[19]);
  CarryOperator U68 (G1[21], P1[21], G0[21], P0[21], G0[20], P0[20]);
  CarryOperator U69 (G1[22], P1[22], G0[22], P0[22], G0[21], P0[21]);
  CarryOperator U70 (G1[23], P1[23], G0[23], P0[23], G0[22], P0[22]);
  CarryOperator U71 (G1[24], P1[24], G0[24], P0[24], G0[23], P0[23]);
  CarryOperator U72 (G1[25], P1[25], G0[25], P0[25], G0[24], P0[24]);
  CarryOperator U73 (G1[26], P1[26], G0[26], P0[26], G0[25], P0[25]);
  CarryOperator U74 (G1[27], P1[27], G0[27], P0[27], G0[26], P0[26]);
  CarryOperator U75 (G1[28], P1[28], G0[28], P0[28], G0[27], P0[27]);
  CarryOperator U76 (G1[29], P1[29], G0[29], P0[29], G0[28], P0[28]);
  CarryOperator U77 (G1[30], P1[30], G0[30], P0[30], G0[29], P0[29]);
  CarryOperator U78 (G1[31], P1[31], G0[31], P0[31], G0[30], P0[30]);
  CarryOperator U79 (G1[32], P1[32], G0[32], P0[32], G0[31], P0[31]);
  CarryOperator U80 (G1[33], P1[33], G0[33], P0[33], G0[32], P0[32]);
  CarryOperator U81 (G1[34], P1[34], G0[34], P0[34], G0[33], P0[33]);
  CarryOperator U82 (G1[35], P1[35], G0[35], P0[35], G0[34], P0[34]);
  CarryOperator U83 (G1[36], P1[36], G0[36], P0[36], G0[35], P0[35]);
  CarryOperator U84 (G1[37], P1[37], G0[37], P0[37], G0[36], P0[36]);
  CarryOperator U85 (G1[38], P1[38], G0[38], P0[38], G0[37], P0[37]);
  CarryOperator U86 (G1[39], P1[39], G0[39], P0[39], G0[38], P0[38]);
  CarryOperator U87 (G1[40], P1[40], G0[40], P0[40], G0[39], P0[39]);
  CarryOperator U88 (G1[41], P1[41], G0[41], P0[41], G0[40], P0[40]);
  CarryOperator U89 (G1[42], P1[42], G0[42], P0[42], G0[41], P0[41]);
  CarryOperator U90 (G1[43], P1[43], G0[43], P0[43], G0[42], P0[42]);
  CarryOperator U91 (G1[44], P1[44], G0[44], P0[44], G0[43], P0[43]);
  CarryOperator U92 (G1[45], P1[45], G0[45], P0[45], G0[44], P0[44]);
  CarryOperator U93 (G1[46], P1[46], G0[46], P0[46], G0[45], P0[45]);
  CarryOperator U94 (G1[47], P1[47], G0[47], P0[47], G0[46], P0[46]);
  CarryOperator U95 (G2[2], P2[2], G1[2], P1[2], G1[0], P1[0]);
  CarryOperator U96 (G2[3], P2[3], G1[3], P1[3], G1[1], P1[1]);
  CarryOperator U97 (G2[4], P2[4], G1[4], P1[4], G1[2], P1[2]);
  CarryOperator U98 (G2[5], P2[5], G1[5], P1[5], G1[3], P1[3]);
  CarryOperator U99 (G2[6], P2[6], G1[6], P1[6], G1[4], P1[4]);
  CarryOperator U100 (G2[7], P2[7], G1[7], P1[7], G1[5], P1[5]);
  CarryOperator U101 (G2[8], P2[8], G1[8], P1[8], G1[6], P1[6]);
  CarryOperator U102 (G2[9], P2[9], G1[9], P1[9], G1[7], P1[7]);
  CarryOperator U103 (G2[10], P2[10], G1[10], P1[10], G1[8], P1[8]);
  CarryOperator U104 (G2[11], P2[11], G1[11], P1[11], G1[9], P1[9]);
  CarryOperator U105 (G2[12], P2[12], G1[12], P1[12], G1[10], P1[10]);
  CarryOperator U106 (G2[13], P2[13], G1[13], P1[13], G1[11], P1[11]);
  CarryOperator U107 (G2[14], P2[14], G1[14], P1[14], G1[12], P1[12]);
  CarryOperator U108 (G2[15], P2[15], G1[15], P1[15], G1[13], P1[13]);
  CarryOperator U109 (G2[16], P2[16], G1[16], P1[16], G1[14], P1[14]);
  CarryOperator U110 (G2[17], P2[17], G1[17], P1[17], G1[15], P1[15]);
  CarryOperator U111 (G2[18], P2[18], G1[18], P1[18], G1[16], P1[16]);
  CarryOperator U112 (G2[19], P2[19], G1[19], P1[19], G1[17], P1[17]);
  CarryOperator U113 (G2[20], P2[20], G1[20], P1[20], G1[18], P1[18]);
  CarryOperator U114 (G2[21], P2[21], G1[21], P1[21], G1[19], P1[19]);
  CarryOperator U115 (G2[22], P2[22], G1[22], P1[22], G1[20], P1[20]);
  CarryOperator U116 (G2[23], P2[23], G1[23], P1[23], G1[21], P1[21]);
  CarryOperator U117 (G2[24], P2[24], G1[24], P1[24], G1[22], P1[22]);
  CarryOperator U118 (G2[25], P2[25], G1[25], P1[25], G1[23], P1[23]);
  CarryOperator U119 (G2[26], P2[26], G1[26], P1[26], G1[24], P1[24]);
  CarryOperator U120 (G2[27], P2[27], G1[27], P1[27], G1[25], P1[25]);
  CarryOperator U121 (G2[28], P2[28], G1[28], P1[28], G1[26], P1[26]);
  CarryOperator U122 (G2[29], P2[29], G1[29], P1[29], G1[27], P1[27]);
  CarryOperator U123 (G2[30], P2[30], G1[30], P1[30], G1[28], P1[28]);
  CarryOperator U124 (G2[31], P2[31], G1[31], P1[31], G1[29], P1[29]);
  CarryOperator U125 (G2[32], P2[32], G1[32], P1[32], G1[30], P1[30]);
  CarryOperator U126 (G2[33], P2[33], G1[33], P1[33], G1[31], P1[31]);
  CarryOperator U127 (G2[34], P2[34], G1[34], P1[34], G1[32], P1[32]);
  CarryOperator U128 (G2[35], P2[35], G1[35], P1[35], G1[33], P1[33]);
  CarryOperator U129 (G2[36], P2[36], G1[36], P1[36], G1[34], P1[34]);
  CarryOperator U130 (G2[37], P2[37], G1[37], P1[37], G1[35], P1[35]);
  CarryOperator U131 (G2[38], P2[38], G1[38], P1[38], G1[36], P1[36]);
  CarryOperator U132 (G2[39], P2[39], G1[39], P1[39], G1[37], P1[37]);
  CarryOperator U133 (G2[40], P2[40], G1[40], P1[40], G1[38], P1[38]);
  CarryOperator U134 (G2[41], P2[41], G1[41], P1[41], G1[39], P1[39]);
  CarryOperator U135 (G2[42], P2[42], G1[42], P1[42], G1[40], P1[40]);
  CarryOperator U136 (G2[43], P2[43], G1[43], P1[43], G1[41], P1[41]);
  CarryOperator U137 (G2[44], P2[44], G1[44], P1[44], G1[42], P1[42]);
  CarryOperator U138 (G2[45], P2[45], G1[45], P1[45], G1[43], P1[43]);
  CarryOperator U139 (G2[46], P2[46], G1[46], P1[46], G1[44], P1[44]);
  CarryOperator U140 (G2[47], P2[47], G1[47], P1[47], G1[45], P1[45]);
  CarryOperator U141 (G3[4], P3[4], G2[4], P2[4], G2[0], P2[0]);
  CarryOperator U142 (G3[5], P3[5], G2[5], P2[5], G2[1], P2[1]);
  CarryOperator U143 (G3[6], P3[6], G2[6], P2[6], G2[2], P2[2]);
  CarryOperator U144 (G3[7], P3[7], G2[7], P2[7], G2[3], P2[3]);
  CarryOperator U145 (G3[8], P3[8], G2[8], P2[8], G2[4], P2[4]);
  CarryOperator U146 (G3[9], P3[9], G2[9], P2[9], G2[5], P2[5]);
  CarryOperator U147 (G3[10], P3[10], G2[10], P2[10], G2[6], P2[6]);
  CarryOperator U148 (G3[11], P3[11], G2[11], P2[11], G2[7], P2[7]);
  CarryOperator U149 (G3[12], P3[12], G2[12], P2[12], G2[8], P2[8]);
  CarryOperator U150 (G3[13], P3[13], G2[13], P2[13], G2[9], P2[9]);
  CarryOperator U151 (G3[14], P3[14], G2[14], P2[14], G2[10], P2[10]);
  CarryOperator U152 (G3[15], P3[15], G2[15], P2[15], G2[11], P2[11]);
  CarryOperator U153 (G3[16], P3[16], G2[16], P2[16], G2[12], P2[12]);
  CarryOperator U154 (G3[17], P3[17], G2[17], P2[17], G2[13], P2[13]);
  CarryOperator U155 (G3[18], P3[18], G2[18], P2[18], G2[14], P2[14]);
  CarryOperator U156 (G3[19], P3[19], G2[19], P2[19], G2[15], P2[15]);
  CarryOperator U157 (G3[20], P3[20], G2[20], P2[20], G2[16], P2[16]);
  CarryOperator U158 (G3[21], P3[21], G2[21], P2[21], G2[17], P2[17]);
  CarryOperator U159 (G3[22], P3[22], G2[22], P2[22], G2[18], P2[18]);
  CarryOperator U160 (G3[23], P3[23], G2[23], P2[23], G2[19], P2[19]);
  CarryOperator U161 (G3[24], P3[24], G2[24], P2[24], G2[20], P2[20]);
  CarryOperator U162 (G3[25], P3[25], G2[25], P2[25], G2[21], P2[21]);
  CarryOperator U163 (G3[26], P3[26], G2[26], P2[26], G2[22], P2[22]);
  CarryOperator U164 (G3[27], P3[27], G2[27], P2[27], G2[23], P2[23]);
  CarryOperator U165 (G3[28], P3[28], G2[28], P2[28], G2[24], P2[24]);
  CarryOperator U166 (G3[29], P3[29], G2[29], P2[29], G2[25], P2[25]);
  CarryOperator U167 (G3[30], P3[30], G2[30], P2[30], G2[26], P2[26]);
  CarryOperator U168 (G3[31], P3[31], G2[31], P2[31], G2[27], P2[27]);
  CarryOperator U169 (G3[32], P3[32], G2[32], P2[32], G2[28], P2[28]);
  CarryOperator U170 (G3[33], P3[33], G2[33], P2[33], G2[29], P2[29]);
  CarryOperator U171 (G3[34], P3[34], G2[34], P2[34], G2[30], P2[30]);
  CarryOperator U172 (G3[35], P3[35], G2[35], P2[35], G2[31], P2[31]);
  CarryOperator U173 (G3[36], P3[36], G2[36], P2[36], G2[32], P2[32]);
  CarryOperator U174 (G3[37], P3[37], G2[37], P2[37], G2[33], P2[33]);
  CarryOperator U175 (G3[38], P3[38], G2[38], P2[38], G2[34], P2[34]);
  CarryOperator U176 (G3[39], P3[39], G2[39], P2[39], G2[35], P2[35]);
  CarryOperator U177 (G3[40], P3[40], G2[40], P2[40], G2[36], P2[36]);
  CarryOperator U178 (G3[41], P3[41], G2[41], P2[41], G2[37], P2[37]);
  CarryOperator U179 (G3[42], P3[42], G2[42], P2[42], G2[38], P2[38]);
  CarryOperator U180 (G3[43], P3[43], G2[43], P2[43], G2[39], P2[39]);
  CarryOperator U181 (G3[44], P3[44], G2[44], P2[44], G2[40], P2[40]);
  CarryOperator U182 (G3[45], P3[45], G2[45], P2[45], G2[41], P2[41]);
  CarryOperator U183 (G3[46], P3[46], G2[46], P2[46], G2[42], P2[42]);
  CarryOperator U184 (G3[47], P3[47], G2[47], P2[47], G2[43], P2[43]);
  CarryOperator U185 (G4[8], P4[8], G3[8], P3[8], G3[0], P3[0]);
  CarryOperator U186 (G4[9], P4[9], G3[9], P3[9], G3[1], P3[1]);
  CarryOperator U187 (G4[10], P4[10], G3[10], P3[10], G3[2], P3[2]);
  CarryOperator U188 (G4[11], P4[11], G3[11], P3[11], G3[3], P3[3]);
  CarryOperator U189 (G4[12], P4[12], G3[12], P3[12], G3[4], P3[4]);
  CarryOperator U190 (G4[13], P4[13], G3[13], P3[13], G3[5], P3[5]);
  CarryOperator U191 (G4[14], P4[14], G3[14], P3[14], G3[6], P3[6]);
  CarryOperator U192 (G4[15], P4[15], G3[15], P3[15], G3[7], P3[7]);
  CarryOperator U193 (G4[16], P4[16], G3[16], P3[16], G3[8], P3[8]);
  CarryOperator U194 (G4[17], P4[17], G3[17], P3[17], G3[9], P3[9]);
  CarryOperator U195 (G4[18], P4[18], G3[18], P3[18], G3[10], P3[10]);
  CarryOperator U196 (G4[19], P4[19], G3[19], P3[19], G3[11], P3[11]);
  CarryOperator U197 (G4[20], P4[20], G3[20], P3[20], G3[12], P3[12]);
  CarryOperator U198 (G4[21], P4[21], G3[21], P3[21], G3[13], P3[13]);
  CarryOperator U199 (G4[22], P4[22], G3[22], P3[22], G3[14], P3[14]);
  CarryOperator U200 (G4[23], P4[23], G3[23], P3[23], G3[15], P3[15]);
  CarryOperator U201 (G4[24], P4[24], G3[24], P3[24], G3[16], P3[16]);
  CarryOperator U202 (G4[25], P4[25], G3[25], P3[25], G3[17], P3[17]);
  CarryOperator U203 (G4[26], P4[26], G3[26], P3[26], G3[18], P3[18]);
  CarryOperator U204 (G4[27], P4[27], G3[27], P3[27], G3[19], P3[19]);
  CarryOperator U205 (G4[28], P4[28], G3[28], P3[28], G3[20], P3[20]);
  CarryOperator U206 (G4[29], P4[29], G3[29], P3[29], G3[21], P3[21]);
  CarryOperator U207 (G4[30], P4[30], G3[30], P3[30], G3[22], P3[22]);
  CarryOperator U208 (G4[31], P4[31], G3[31], P3[31], G3[23], P3[23]);
  CarryOperator U209 (G4[32], P4[32], G3[32], P3[32], G3[24], P3[24]);
  CarryOperator U210 (G4[33], P4[33], G3[33], P3[33], G3[25], P3[25]);
  CarryOperator U211 (G4[34], P4[34], G3[34], P3[34], G3[26], P3[26]);
  CarryOperator U212 (G4[35], P4[35], G3[35], P3[35], G3[27], P3[27]);
  CarryOperator U213 (G4[36], P4[36], G3[36], P3[36], G3[28], P3[28]);
  CarryOperator U214 (G4[37], P4[37], G3[37], P3[37], G3[29], P3[29]);
  CarryOperator U215 (G4[38], P4[38], G3[38], P3[38], G3[30], P3[30]);
  CarryOperator U216 (G4[39], P4[39], G3[39], P3[39], G3[31], P3[31]);
  CarryOperator U217 (G4[40], P4[40], G3[40], P3[40], G3[32], P3[32]);
  CarryOperator U218 (G4[41], P4[41], G3[41], P3[41], G3[33], P3[33]);
  CarryOperator U219 (G4[42], P4[42], G3[42], P3[42], G3[34], P3[34]);
  CarryOperator U220 (G4[43], P4[43], G3[43], P3[43], G3[35], P3[35]);
  CarryOperator U221 (G4[44], P4[44], G3[44], P3[44], G3[36], P3[36]);
  CarryOperator U222 (G4[45], P4[45], G3[45], P3[45], G3[37], P3[37]);
  CarryOperator U223 (G4[46], P4[46], G3[46], P3[46], G3[38], P3[38]);
  CarryOperator U224 (G4[47], P4[47], G3[47], P3[47], G3[39], P3[39]);
  CarryOperator U225 (G5[16], P5[16], G4[16], P4[16], G4[0], P4[0]);
  CarryOperator U226 (G5[17], P5[17], G4[17], P4[17], G4[1], P4[1]);
  CarryOperator U227 (G5[18], P5[18], G4[18], P4[18], G4[2], P4[2]);
  CarryOperator U228 (G5[19], P5[19], G4[19], P4[19], G4[3], P4[3]);
  CarryOperator U229 (G5[20], P5[20], G4[20], P4[20], G4[4], P4[4]);
  CarryOperator U230 (G5[21], P5[21], G4[21], P4[21], G4[5], P4[5]);
  CarryOperator U231 (G5[22], P5[22], G4[22], P4[22], G4[6], P4[6]);
  CarryOperator U232 (G5[23], P5[23], G4[23], P4[23], G4[7], P4[7]);
  CarryOperator U233 (G5[24], P5[24], G4[24], P4[24], G4[8], P4[8]);
  CarryOperator U234 (G5[25], P5[25], G4[25], P4[25], G4[9], P4[9]);
  CarryOperator U235 (G5[26], P5[26], G4[26], P4[26], G4[10], P4[10]);
  CarryOperator U236 (G5[27], P5[27], G4[27], P4[27], G4[11], P4[11]);
  CarryOperator U237 (G5[28], P5[28], G4[28], P4[28], G4[12], P4[12]);
  CarryOperator U238 (G5[29], P5[29], G4[29], P4[29], G4[13], P4[13]);
  CarryOperator U239 (G5[30], P5[30], G4[30], P4[30], G4[14], P4[14]);
  CarryOperator U240 (G5[31], P5[31], G4[31], P4[31], G4[15], P4[15]);
  CarryOperator U241 (G5[32], P5[32], G4[32], P4[32], G4[16], P4[16]);
  CarryOperator U242 (G5[33], P5[33], G4[33], P4[33], G4[17], P4[17]);
  CarryOperator U243 (G5[34], P5[34], G4[34], P4[34], G4[18], P4[18]);
  CarryOperator U244 (G5[35], P5[35], G4[35], P4[35], G4[19], P4[19]);
  CarryOperator U245 (G5[36], P5[36], G4[36], P4[36], G4[20], P4[20]);
  CarryOperator U246 (G5[37], P5[37], G4[37], P4[37], G4[21], P4[21]);
  CarryOperator U247 (G5[38], P5[38], G4[38], P4[38], G4[22], P4[22]);
  CarryOperator U248 (G5[39], P5[39], G4[39], P4[39], G4[23], P4[23]);
  CarryOperator U249 (G5[40], P5[40], G4[40], P4[40], G4[24], P4[24]);
  CarryOperator U250 (G5[41], P5[41], G4[41], P4[41], G4[25], P4[25]);
  CarryOperator U251 (G5[42], P5[42], G4[42], P4[42], G4[26], P4[26]);
  CarryOperator U252 (G5[43], P5[43], G4[43], P4[43], G4[27], P4[27]);
  CarryOperator U253 (G5[44], P5[44], G4[44], P4[44], G4[28], P4[28]);
  CarryOperator U254 (G5[45], P5[45], G4[45], P4[45], G4[29], P4[29]);
  CarryOperator U255 (G5[46], P5[46], G4[46], P4[46], G4[30], P4[30]);
  CarryOperator U256 (G5[47], P5[47], G4[47], P4[47], G4[31], P4[31]);
  CarryOperator U257 (G6[32], P6[32], G5[32], P5[32], G5[0], P5[0]);
  CarryOperator U258 (G6[33], P6[33], G5[33], P5[33], G5[1], P5[1]);
  CarryOperator U259 (G6[34], P6[34], G5[34], P5[34], G5[2], P5[2]);
  CarryOperator U260 (G6[35], P6[35], G5[35], P5[35], G5[3], P5[3]);
  CarryOperator U261 (G6[36], P6[36], G5[36], P5[36], G5[4], P5[4]);
  CarryOperator U262 (G6[37], P6[37], G5[37], P5[37], G5[5], P5[5]);
  CarryOperator U263 (G6[38], P6[38], G5[38], P5[38], G5[6], P5[6]);
  CarryOperator U264 (G6[39], P6[39], G5[39], P5[39], G5[7], P5[7]);
  CarryOperator U265 (G6[40], P6[40], G5[40], P5[40], G5[8], P5[8]);
  CarryOperator U266 (G6[41], P6[41], G5[41], P5[41], G5[9], P5[9]);
  CarryOperator U267 (G6[42], P6[42], G5[42], P5[42], G5[10], P5[10]);
  CarryOperator U268 (G6[43], P6[43], G5[43], P5[43], G5[11], P5[11]);
  CarryOperator U269 (G6[44], P6[44], G5[44], P5[44], G5[12], P5[12]);
  CarryOperator U270 (G6[45], P6[45], G5[45], P5[45], G5[13], P5[13]);
  CarryOperator U271 (G6[46], P6[46], G5[46], P5[46], G5[14], P5[14]);
  CarryOperator U272 (G6[47], P6[47], G5[47], P5[47], G5[15], P5[15]);
endmodule

module UBZero_0_0(O);
  output [0:0] O;
  assign O[0] = 0;
endmodule

module UBCON_31_0 (O, I);
  output [31:0] O;
  input [31:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
  UB1DCON_13 U13 (O[13], I[13]);
  UB1DCON_14 U14 (O[14], I[14]);
  UB1DCON_15 U15 (O[15], I[15]);
  UB1DCON_16 U16 (O[16], I[16]);
  UB1DCON_17 U17 (O[17], I[17]);
  UB1DCON_18 U18 (O[18], I[18]);
  UB1DCON_19 U19 (O[19], I[19]);
  UB1DCON_20 U20 (O[20], I[20]);
  UB1DCON_21 U21 (O[21], I[21]);
  UB1DCON_22 U22 (O[22], I[22]);
  UB1DCON_23 U23 (O[23], I[23]);
  UB1DCON_24 U24 (O[24], I[24]);
  UB1DCON_25 U25 (O[25], I[25]);
  UB1DCON_26 U26 (O[26], I[26]);
  UB1DCON_27 U27 (O[27], I[27]);
  UB1DCON_28 U28 (O[28], I[28]);
  UB1DCON_29 U29 (O[29], I[29]);
  UB1DCON_30 U30 (O[30], I[30]);
  UB1DCON_31 U31 (O[31], I[31]);
endmodule

module UBExtender_31_0_4000 (O, I);
  output [47:0] O;
  input [31:0] I;
  UBCON_31_0 U0 (O[31:0], I[31:0]);
  UBZero_47_32 U1 (O[47:32]);
endmodule

module UBKSA_31_0_47_0 (S, X, Y);
  output [48:0] S;
  input [31:0] X;
  input [47:0] Y;
  wire [47:0] Z;
  UBExtender_31_0_4000 U0 (Z[47:0], X[31:0]);
  UBPureKSA_47_0 U1 (S[48:0], Z[47:0], Y[47:0]);
endmodule

module UBPureKSA_47_0 (S, X, Y);
  output [48:0] S;
  input [47:0] X;
  input [47:0] Y;
  wire C;
  UBPriKSA_47_0 U0 (S, X, Y, C);
  UBZero_0_0 U1 (C);
endmodule

