/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: Multiplier_15_0_1000

  Number system: Unsigned binary
  Multiplicand length: 16
  Multiplier length: 16
  Partial product generation: Simple PPG
  Partial product accumulation: Overturned-stairs tree
  Final stage addition: Carry-skip adder (fixed-block-size)
----------------------------------------------------------------------------*/

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_1(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_2(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_12(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_13(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_14(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_15(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_16(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_16(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_17(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_18(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_19(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_7(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_19(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_20(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_21(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_22(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_23(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_6(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_21(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_23(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_5(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_20(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_21(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_24(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_10(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_22(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_23(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_24(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_25(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_11(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_25(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_26(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB1DCON_27(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_9(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_24(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_26(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_27(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_8(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_25(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_28(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_14(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_27(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_28(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_29(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_30(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_13(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_28(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_30(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_12(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_29(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_31(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBFA_29(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBPFA_4(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_4 U0 (C_0, S_0, X, Y);
  UBHA_4 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_5(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_5 U0 (C_0, S_0, X, Y);
  UBHA_5 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_6(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_6 U0 (C_0, S_0, X, Y);
  UBHA_6 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_6_4(Co, S, X, Y, Ci);
  output Co;
  output [6:4] S;
  input Ci;
  input [6:4] X;
  input [6:4] Y;
  wire C5;
  wire C6;
  wire C7;
  wire P4;
  wire P5;
  wire P6;
  wire Sk;
  assign Sk = ( P4 & P5 & P6 ) & Ci;
  assign Co = C7 | Sk;
  UBPFA_4 U0 (C5, S[4], P4, X[4], Y[4], Ci);
  UBPFA_5 U1 (C6, S[5], P5, X[5], Y[5], C5);
  UBPFA_6 U2 (C7, S[6], P6, X[6], Y[6], C6);
endmodule

module UBPFA_7(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_7 U0 (C_0, S_0, X, Y);
  UBHA_7 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_8(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_8 U0 (C_0, S_0, X, Y);
  UBHA_8 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_9(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_9 U0 (C_0, S_0, X, Y);
  UBHA_9 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_9_7(Co, S, X, Y, Ci);
  output Co;
  output [9:7] S;
  input Ci;
  input [9:7] X;
  input [9:7] Y;
  wire C10;
  wire C8;
  wire C9;
  wire P7;
  wire P8;
  wire P9;
  wire Sk;
  assign Sk = ( P7 & P8 & P9 ) & Ci;
  assign Co = C10 | Sk;
  UBPFA_7 U0 (C8, S[7], P7, X[7], Y[7], Ci);
  UBPFA_8 U1 (C9, S[8], P8, X[8], Y[8], C8);
  UBPFA_9 U2 (C10, S[9], P9, X[9], Y[9], C9);
endmodule

module UBPFA_10(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_10 U0 (C_0, S_0, X, Y);
  UBHA_10 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_11(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_11 U0 (C_0, S_0, X, Y);
  UBHA_11 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_12(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_12 U0 (C_0, S_0, X, Y);
  UBHA_12 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_12_10(Co, S, X, Y, Ci);
  output Co;
  output [12:10] S;
  input Ci;
  input [12:10] X;
  input [12:10] Y;
  wire C11;
  wire C12;
  wire C13;
  wire P10;
  wire P11;
  wire P12;
  wire Sk;
  assign Sk = ( P10 & P11 & P12 ) & Ci;
  assign Co = C13 | Sk;
  UBPFA_10 U0 (C11, S[10], P10, X[10], Y[10], Ci);
  UBPFA_11 U1 (C12, S[11], P11, X[11], Y[11], C11);
  UBPFA_12 U2 (C13, S[12], P12, X[12], Y[12], C12);
endmodule

module UBPFA_13(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_13 U0 (C_0, S_0, X, Y);
  UBHA_13 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_14(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_14 U0 (C_0, S_0, X, Y);
  UBHA_14 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_15(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_15(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_15 U0 (C_0, S_0, X, Y);
  UBHA_15 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_15_13(Co, S, X, Y, Ci);
  output Co;
  output [15:13] S;
  input Ci;
  input [15:13] X;
  input [15:13] Y;
  wire C14;
  wire C15;
  wire C16;
  wire P13;
  wire P14;
  wire P15;
  wire Sk;
  assign Sk = ( P13 & P14 & P15 ) & Ci;
  assign Co = C16 | Sk;
  UBPFA_13 U0 (C14, S[13], P13, X[13], Y[13], Ci);
  UBPFA_14 U1 (C15, S[14], P14, X[14], Y[14], C14);
  UBPFA_15 U2 (C16, S[15], P15, X[15], Y[15], C15);
endmodule

module UBPFA_16(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_16 U0 (C_0, S_0, X, Y);
  UBHA_16 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_17(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_17(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_17 U0 (C_0, S_0, X, Y);
  UBHA_17 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_18(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_18(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_18 U0 (C_0, S_0, X, Y);
  UBHA_18 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_18_16(Co, S, X, Y, Ci);
  output Co;
  output [18:16] S;
  input Ci;
  input [18:16] X;
  input [18:16] Y;
  wire C17;
  wire C18;
  wire C19;
  wire P16;
  wire P17;
  wire P18;
  wire Sk;
  assign Sk = ( P16 & P17 & P18 ) & Ci;
  assign Co = C19 | Sk;
  UBPFA_16 U0 (C17, S[16], P16, X[16], Y[16], Ci);
  UBPFA_17 U1 (C18, S[17], P17, X[17], Y[17], C17);
  UBPFA_18 U2 (C19, S[18], P18, X[18], Y[18], C18);
endmodule

module UBPFA_19(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_19 U0 (C_0, S_0, X, Y);
  UBHA_19 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_20(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_20 U0 (C_0, S_0, X, Y);
  UBHA_20 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_21(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_21 U0 (C_0, S_0, X, Y);
  UBHA_21 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_21_19(Co, S, X, Y, Ci);
  output Co;
  output [21:19] S;
  input Ci;
  input [21:19] X;
  input [21:19] Y;
  wire C20;
  wire C21;
  wire C22;
  wire P19;
  wire P20;
  wire P21;
  wire Sk;
  assign Sk = ( P19 & P20 & P21 ) & Ci;
  assign Co = C22 | Sk;
  UBPFA_19 U0 (C20, S[19], P19, X[19], Y[19], Ci);
  UBPFA_20 U1 (C21, S[20], P20, X[20], Y[20], C20);
  UBPFA_21 U2 (C22, S[21], P21, X[21], Y[21], C21);
endmodule

module UBPFA_22(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_22 U0 (C_0, S_0, X, Y);
  UBHA_22 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_23(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_23 U0 (C_0, S_0, X, Y);
  UBHA_23 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_24(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_24 U0 (C_0, S_0, X, Y);
  UBHA_24 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_24_22(Co, S, X, Y, Ci);
  output Co;
  output [24:22] S;
  input Ci;
  input [24:22] X;
  input [24:22] Y;
  wire C23;
  wire C24;
  wire C25;
  wire P22;
  wire P23;
  wire P24;
  wire Sk;
  assign Sk = ( P22 & P23 & P24 ) & Ci;
  assign Co = C25 | Sk;
  UBPFA_22 U0 (C23, S[22], P22, X[22], Y[22], Ci);
  UBPFA_23 U1 (C24, S[23], P23, X[23], Y[23], C23);
  UBPFA_24 U2 (C25, S[24], P24, X[24], Y[24], C24);
endmodule

module UBPFA_25(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_25 U0 (C_0, S_0, X, Y);
  UBHA_25 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_26(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_26 U0 (C_0, S_0, X, Y);
  UBHA_26 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_27(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_27 U0 (C_0, S_0, X, Y);
  UBHA_27 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_27_25(Co, S, X, Y, Ci);
  output Co;
  output [27:25] S;
  input Ci;
  input [27:25] X;
  input [27:25] Y;
  wire C26;
  wire C27;
  wire C28;
  wire P25;
  wire P26;
  wire P27;
  wire Sk;
  assign Sk = ( P25 & P26 & P27 ) & Ci;
  assign Co = C28 | Sk;
  UBPFA_25 U0 (C26, S[25], P25, X[25], Y[25], Ci);
  UBPFA_26 U1 (C27, S[26], P26, X[26], Y[26], C26);
  UBPFA_27 U2 (C28, S[27], P27, X[27], Y[27], C27);
endmodule

module UBPFA_28(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_28 U0 (C_0, S_0, X, Y);
  UBHA_28 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_29(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_29 U0 (C_0, S_0, X, Y);
  UBHA_29 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_30(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_30 U0 (C_0, S_0, X, Y);
  UBHA_30 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_30_28(Co, S, X, Y, Ci);
  output Co;
  output [30:28] S;
  input Ci;
  input [30:28] X;
  input [30:28] Y;
  wire C29;
  wire C30;
  wire C31;
  wire P28;
  wire P29;
  wire P30;
  wire Sk;
  assign Sk = ( P28 & P29 & P30 ) & Ci;
  assign Co = C31 | Sk;
  UBPFA_28 U0 (C29, S[28], P28, X[28], Y[28], Ci);
  UBPFA_29 U1 (C30, S[29], P29, X[29], Y[29], C29);
  UBPFA_30 U2 (C31, S[30], P30, X[30], Y[30], C30);
endmodule

module UBHA_31(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_31(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_31 U0 (C_0, S_0, X, Y);
  UBHA_31 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_31_31(Co, S, X, Y, Ci);
  output Co;
  output [31:31] S;
  input Ci;
  input [31:31] X;
  input [31:31] Y;
  wire C32;
  wire P31;
  wire Sk;
  assign Sk = P31 & Ci;
  assign Co = C32 | Sk;
  UBPFA_31 U0 (C32, S[31], P31, X[31], Y[31], Ci);
endmodule

module UBPriFCSkA_31_4(S, X, Y, Cin);
  output [32:4] S;
  input Cin;
  input [31:4] X;
  input [31:4] Y;
  wire C10;
  wire C13;
  wire C16;
  wire C19;
  wire C22;
  wire C25;
  wire C28;
  wire C31;
  wire C7;
  UBCSkB_6_4 U0 (C7, S[6:4], X[6:4], Y[6:4], Cin);
  UBCSkB_9_7 U1 (C10, S[9:7], X[9:7], Y[9:7], C7);
  UBCSkB_12_10 U2 (C13, S[12:10], X[12:10], Y[12:10], C10);
  UBCSkB_15_13 U3 (C16, S[15:13], X[15:13], Y[15:13], C13);
  UBCSkB_18_16 U4 (C19, S[18:16], X[18:16], Y[18:16], C16);
  UBCSkB_21_19 U5 (C22, S[21:19], X[21:19], Y[21:19], C19);
  UBCSkB_24_22 U6 (C25, S[24:22], X[24:22], Y[24:22], C22);
  UBCSkB_27_25 U7 (C28, S[27:25], X[27:25], Y[27:25], C25);
  UBCSkB_30_28 U8 (C31, S[30:28], X[30:28], Y[30:28], C28);
  UBCSkB_31_31 U9 (S[32], S[31], X[31], Y[31], C31);
endmodule

module UBZero_4_4(O);
  output [4:4] O;
  assign O[4] = 0;
endmodule

module Multiplier_15_0_1000(P, IN1, IN2);
  output [31:0] P;
  input [15:0] IN1;
  input [15:0] IN2;
  wire [32:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  assign P[12] = W[12];
  assign P[13] = W[13];
  assign P[14] = W[14];
  assign P[15] = W[15];
  assign P[16] = W[16];
  assign P[17] = W[17];
  assign P[18] = W[18];
  assign P[19] = W[19];
  assign P[20] = W[20];
  assign P[21] = W[21];
  assign P[22] = W[22];
  assign P[23] = W[23];
  assign P[24] = W[24];
  assign P[25] = W[25];
  assign P[26] = W[26];
  assign P[27] = W[27];
  assign P[28] = W[28];
  assign P[29] = W[29];
  assign P[30] = W[30];
  assign P[31] = W[31];
  MultUB_STD_OS_FCS000 U0 (W, IN1, IN2);
endmodule

module CSA_15_0_16_1_17_000 (C, S, X, Y, Z);
  output [17:2] C;
  output [17:0] S;
  input [15:0] X;
  input [16:1] Y;
  input [17:2] Z;
  UB1DCON_0 U0 (S[0], X[0]);
  UBHA_1 U1 (C[2], S[1], Y[1], X[1]);
  PureCSA_15_2 U2 (C[16:3], S[15:2], Z[15:2], Y[15:2], X[15:2]);
  UBHA_16 U3 (C[17], S[16], Z[16], Y[16]);
  UB1DCON_17 U4 (S[17], Z[17]);
endmodule

module CSA_17_2_17_0_20_000 (C, S, X, Y, Z);
  output [18:3] C;
  output [20:0] S;
  input [17:2] X;
  input [17:0] Y;
  input [20:5] Z;
  UBCON_1_0 U0 (S[1:0], Y[1:0]);
  PureCSHA_4_2 U1 (C[5:3], S[4:2], X[4:2], Y[4:2]);
  PureCSA_17_5 U2 (C[18:6], S[17:5], Z[17:5], X[17:5], Y[17:5]);
  UBCON_20_18 U3 (S[20:18], Z[20:18]);
endmodule

module CSA_18_3_19_4_20_000 (C, S, X, Y, Z);
  output [20:5] C;
  output [20:3] S;
  input [18:3] X;
  input [19:4] Y;
  input [20:5] Z;
  UB1DCON_3 U0 (S[3], X[3]);
  UBHA_4 U1 (C[5], S[4], Y[4], X[4]);
  PureCSA_18_5 U2 (C[19:6], S[18:5], Z[18:5], Y[18:5], X[18:5]);
  UBHA_19 U3 (C[20], S[19], Z[19], Y[19]);
  UB1DCON_20 U4 (S[20], Z[20]);
endmodule

module CSA_18_3_20_0_24_000 (C, S, X, Y, Z);
  output [21:4] C;
  output [24:0] S;
  input [18:3] X;
  input [20:0] Y;
  input [24:7] Z;
  UBCON_2_0 U0 (S[2:0], Y[2:0]);
  PureCSHA_6_3 U1 (C[7:4], S[6:3], X[6:3], Y[6:3]);
  PureCSA_18_7 U2 (C[19:8], S[18:7], Z[18:7], X[18:7], Y[18:7]);
  PureCSHA_20_19 U3 (C[21:20], S[20:19], Z[20:19], Y[20:19]);
  UBCON_24_21 U4 (S[24:21], Z[24:21]);
endmodule

module CSA_20_3_23_8_23_000 (C, S, X, Y, Z);
  output [24:7] C;
  output [23:3] S;
  input [20:3] X;
  input [23:8] Y;
  input [23:6] Z;
  UBCON_5_3 U0 (S[5:3], X[5:3]);
  PureCSHA_7_6 U1 (C[8:7], S[7:6], Z[7:6], X[7:6]);
  PureCSA_20_8 U2 (C[21:9], S[20:8], Y[20:8], Z[20:8], X[20:8]);
  PureCSHA_23_21 U3 (C[24:22], S[23:21], Z[23:21], Y[23:21]);
endmodule

module CSA_21_4_24_0_28_000 (C, S, X, Y, Z);
  output [25:5] C;
  output [28:0] S;
  input [21:4] X;
  input [24:0] Y;
  input [28:10] Z;
  UBCON_3_0 U0 (S[3:0], Y[3:0]);
  PureCSHA_9_4 U1 (C[10:5], S[9:4], X[9:4], Y[9:4]);
  PureCSA_21_10 U2 (C[22:11], S[21:10], Z[21:10], X[21:10], Y[21:10]);
  PureCSHA_24_22 U3 (C[25:23], S[24:22], Z[24:22], Y[24:22]);
  UBCON_28_25 U4 (S[28:25], Z[28:25]);
endmodule

module CSA_21_6_22_7_23_000 (C, S, X, Y, Z);
  output [23:8] C;
  output [23:6] S;
  input [21:6] X;
  input [22:7] Y;
  input [23:8] Z;
  UB1DCON_6 U0 (S[6], X[6]);
  UBHA_7 U1 (C[8], S[7], Y[7], X[7]);
  PureCSA_21_8 U2 (C[22:9], S[21:8], Z[21:8], Y[21:8], X[21:8]);
  UBHA_22 U3 (C[23], S[22], Z[22], Y[22]);
  UB1DCON_23 U4 (S[23], Z[23]);
endmodule

module CSA_23_3_27_12_27000 (C, S, X, Y, Z);
  output [28:10] C;
  output [27:3] S;
  input [23:3] X;
  input [27:12] Y;
  input [27:9] Z;
  UBCON_8_3 U0 (S[8:3], X[8:3]);
  PureCSHA_11_9 U1 (C[12:10], S[11:9], Z[11:9], X[11:9]);
  PureCSA_23_12 U2 (C[24:13], S[23:12], Y[23:12], Z[23:12], X[23:12]);
  PureCSHA_27_24 U3 (C[28:25], S[27:24], Z[27:24], Y[27:24]);
endmodule

module CSA_24_9_25_10_26000 (C, S, X, Y, Z);
  output [26:11] C;
  output [26:9] S;
  input [24:9] X;
  input [25:10] Y;
  input [26:11] Z;
  UB1DCON_9 U0 (S[9], X[9]);
  UBHA_10 U1 (C[11], S[10], Y[10], X[10]);
  PureCSA_24_11 U2 (C[25:12], S[24:11], Z[24:11], Y[24:11], X[24:11]);
  UBHA_25 U3 (C[26], S[25], Z[25], Y[25]);
  UB1DCON_26 U4 (S[26], Z[26]);
endmodule

module CSA_25_5_28_0_31_000 (C, S, X, Y, Z);
  output [29:6] C;
  output [31:0] S;
  input [25:5] X;
  input [28:0] Y;
  input [31:14] Z;
  UBCON_4_0 U0 (S[4:0], Y[4:0]);
  PureCSHA_13_5 U1 (C[14:6], S[13:5], X[13:5], Y[13:5]);
  PureCSA_25_14 U2 (C[26:15], S[25:14], Z[25:14], X[25:14], Y[25:14]);
  PureCSHA_28_26 U3 (C[29:27], S[28:26], Z[28:26], Y[28:26]);
  UBCON_31_29 U4 (S[31:29], Z[31:29]);
endmodule

module CSA_26_9_26_11_27000 (C, S, X, Y, Z);
  output [27:12] C;
  output [27:9] S;
  input [26:9] X;
  input [26:11] Y;
  input [27:12] Z;
  UBCON_10_9 U0 (S[10:9], X[10:9]);
  UBHA_11 U1 (C[12], S[11], Y[11], X[11]);
  PureCSA_26_12 U2 (C[27:13], S[26:12], Z[26:12], Y[26:12], X[26:12]);
  UB1DCON_27 U3 (S[27], Z[27]);
endmodule

module CSA_27_3_30_15_30000 (C, S, X, Y, Z);
  output [31:14] C;
  output [30:3] S;
  input [27:3] X;
  input [30:15] Y;
  input [30:13] Z;
  UBCON_12_3 U0 (S[12:3], X[12:3]);
  PureCSHA_14_13 U1 (C[15:14], S[14:13], Z[14:13], X[14:13]);
  PureCSA_27_15 U2 (C[28:16], S[27:15], Y[27:15], Z[27:15], X[27:15]);
  PureCSHA_30_28 U3 (C[31:29], S[30:28], Z[30:28], Y[30:28]);
endmodule

module CSA_28_13_29_14_3000 (C, S, X, Y, Z);
  output [30:15] C;
  output [30:13] S;
  input [28:13] X;
  input [29:14] Y;
  input [30:15] Z;
  UB1DCON_13 U0 (S[13], X[13]);
  UBHA_14 U1 (C[15], S[14], Y[14], X[14]);
  PureCSA_28_15 U2 (C[29:16], S[28:15], Z[28:15], Y[28:15], X[28:15]);
  UBHA_29 U3 (C[30], S[29], Z[29], Y[29]);
  UB1DCON_30 U4 (S[30], Z[30]);
endmodule

module CSA_29_6_31_0_30_000 (C, S, X, Y, Z);
  output [31:4] C;
  output [31:0] S;
  input [29:6] X;
  input [31:0] Y;
  input [30:3] Z;
  UBCON_2_0 U0 (S[2:0], Y[2:0]);
  PureCSHA_5_3 U1 (C[6:4], S[5:3], Z[5:3], Y[5:3]);
  PureCSA_29_6 U2 (C[30:7], S[29:6], X[29:6], Z[29:6], Y[29:6]);
  UBHA_30 U3 (C[31], S[30], Y[30], Z[30]);
  UB1DCON_31 U4 (S[31], Y[31]);
endmodule

module MultUB_STD_OS_FCS000 (P, IN1, IN2);
  output [32:0] P;
  input [15:0] IN1;
  input [15:0] IN2;
  wire [15:0] PP0;
  wire [16:1] PP1;
  wire [25:10] PP10;
  wire [26:11] PP11;
  wire [27:12] PP12;
  wire [28:13] PP13;
  wire [29:14] PP14;
  wire [30:15] PP15;
  wire [17:2] PP2;
  wire [18:3] PP3;
  wire [19:4] PP4;
  wire [20:5] PP5;
  wire [21:6] PP6;
  wire [22:7] PP7;
  wire [23:8] PP8;
  wire [24:9] PP9;
  wire [31:4] S1;
  wire [31:0] S2;
  UBPPG_15_0_15_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, IN1, IN2);
  OSTR_15_0_16_1_17000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15);
  UBFCSkA_31_4_31_0 U2 (P, S1, S2);
endmodule

module OSBODY_15_0_16_1_000 (S0, S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15);
  output [29:6] S0;
  output [31:0] S1;
  output [30:3] S2;
  input [15:0] PP0;
  input [16:1] PP1;
  input [25:10] PP10;
  input [26:11] PP11;
  input [27:12] PP12;
  input [28:13] PP13;
  input [29:14] PP14;
  input [30:15] PP15;
  input [17:2] PP2;
  input [18:3] PP3;
  input [19:4] PP4;
  input [20:5] PP5;
  input [21:6] PP6;
  input [22:7] PP7;
  input [23:8] PP8;
  input [24:9] PP9;
  wire [25:5] W0;
  wire [28:0] W1;
  wire [27:3] W2;
  wire [30:15] W3;
  wire [30:13] W4;
  OSBODY_15_0_16_1_001 U0 (W0, W1, W2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12);
  UBARYACC_28_13_29000 U1 (W3, W4, PP13, PP14, PP15);
  OSCON_25_5_28_0_2000 U2 (S0, S1, S2, W0, W1, W2, W3, W4);
endmodule

module OSBODY_15_0_16_1_001 (S0, S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12);
  output [25:5] S0;
  output [28:0] S1;
  output [27:3] S2;
  input [15:0] PP0;
  input [16:1] PP1;
  input [25:10] PP10;
  input [26:11] PP11;
  input [27:12] PP12;
  input [17:2] PP2;
  input [18:3] PP3;
  input [19:4] PP4;
  input [20:5] PP5;
  input [21:6] PP6;
  input [22:7] PP7;
  input [23:8] PP8;
  input [24:9] PP9;
  wire [21:4] W0;
  wire [24:0] W1;
  wire [23:3] W2;
  wire [27:12] W3;
  wire [27:9] W4;
  OSBODY_15_0_16_1_002 U0 (W0, W1, W2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8);
  UBARYACC_24_9_25_000 U1 (W3, W4, PP9, PP10, PP11, PP12);
  OSCON_21_4_24_0_2000 U2 (S0, S1, S2, W0, W1, W2, W3, W4);
endmodule

module OSBODY_15_0_16_1_002 (S0, S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8);
  output [21:4] S0;
  output [24:0] S1;
  output [23:3] S2;
  input [15:0] PP0;
  input [16:1] PP1;
  input [17:2] PP2;
  input [18:3] PP3;
  input [19:4] PP4;
  input [20:5] PP5;
  input [21:6] PP6;
  input [22:7] PP7;
  input [23:8] PP8;
  wire [18:3] W0;
  wire [20:0] W1;
  wire [20:3] W2;
  wire [23:8] W3;
  wire [23:6] W4;
  OSBODY_15_0_16_1_003 U0 (W0, W1, W2, PP0, PP1, PP2, PP3, PP4, PP5);
  UBARYACC_21_6_22_000 U1 (W3, W4, PP6, PP7, PP8);
  OSCON_18_3_20_0_2000 U2 (S0, S1, S2, W0, W1, W2, W3, W4);
endmodule

module OSBODY_15_0_16_1_003 (S0, S1, S2, PP0, PP1, PP2, PP3, PP4, PP5);
  output [18:3] S0;
  output [20:0] S1;
  output [20:3] S2;
  input [15:0] PP0;
  input [16:1] PP1;
  input [17:2] PP2;
  input [18:3] PP3;
  input [19:4] PP4;
  input [20:5] PP5;
  wire [17:2] W0;
  wire [17:0] W1;
  wire [18:3] W2;
  wire [19:4] W3;
  wire [20:5] W4;
  OSBODY_15_0_16_1_004 U0 (W0, W1, W2, PP0, PP1, PP2, PP3);
  UBARYACC_19_4_20_000 U1 (W3, W4, PP4, PP5);
  OSCON_17_2_17_0_1000 U2 (S0, S1, S2, W0, W1, W2, W3, W4);
endmodule

module OSBODY_15_0_16_1_004 (S0, S1, S2, PP0, PP1, PP2, PP3);
  output [17:2] S0;
  output [17:0] S1;
  output [18:3] S2;
  input [15:0] PP0;
  input [16:1] PP1;
  input [17:2] PP2;
  input [18:3] PP3;
  CSA_15_0_16_1_17_000 U0 (S0, S1, PP0, PP1, PP2);
  UBCON_18_3 U1 (S2, PP3);
endmodule

module OSCON_17_2_17_0_1000 (S0, S1, S2, IN0, IN1, IN2, IN3, IN4);
  output [18:3] S0;
  output [20:0] S1;
  output [20:3] S2;
  input [17:2] IN0;
  input [17:0] IN1;
  input [18:3] IN2;
  input [19:4] IN3;
  input [20:5] IN4;
  wire [20:5] W;
  CSA_18_3_19_4_20_000 U0 (W, S2, IN2, IN3, IN4);
  CSA_17_2_17_0_20_000 U1 (S0, S1, IN0, IN1, W);
endmodule

module OSCON_18_3_20_0_2000 (S0, S1, S2, IN0, IN1, IN2, IN3, IN4);
  output [21:4] S0;
  output [24:0] S1;
  output [23:3] S2;
  input [18:3] IN0;
  input [20:0] IN1;
  input [20:3] IN2;
  input [23:8] IN3;
  input [23:6] IN4;
  wire [24:7] W;
  CSA_20_3_23_8_23_000 U0 (W, S2, IN2, IN3, IN4);
  CSA_18_3_20_0_24_000 U1 (S0, S1, IN0, IN1, W);
endmodule

module OSCON_21_4_24_0_2000 (S0, S1, S2, IN0, IN1, IN2, IN3, IN4);
  output [25:5] S0;
  output [28:0] S1;
  output [27:3] S2;
  input [21:4] IN0;
  input [24:0] IN1;
  input [23:3] IN2;
  input [27:12] IN3;
  input [27:9] IN4;
  wire [28:10] W;
  CSA_23_3_27_12_27000 U0 (W, S2, IN2, IN3, IN4);
  CSA_21_4_24_0_28_000 U1 (S0, S1, IN0, IN1, W);
endmodule

module OSCON_25_5_28_0_2000 (S0, S1, S2, IN0, IN1, IN2, IN3, IN4);
  output [29:6] S0;
  output [31:0] S1;
  output [30:3] S2;
  input [25:5] IN0;
  input [28:0] IN1;
  input [27:3] IN2;
  input [30:15] IN3;
  input [30:13] IN4;
  wire [31:14] W;
  CSA_27_3_30_15_30000 U0 (W, S2, IN2, IN3, IN4);
  CSA_25_5_28_0_31_000 U1 (S0, S1, IN0, IN1, W);
endmodule

module OSTR_15_0_16_1_17000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15);
  output [31:4] S1;
  output [31:0] S2;
  input [15:0] PP0;
  input [16:1] PP1;
  input [25:10] PP10;
  input [26:11] PP11;
  input [27:12] PP12;
  input [28:13] PP13;
  input [29:14] PP14;
  input [30:15] PP15;
  input [17:2] PP2;
  input [18:3] PP3;
  input [19:4] PP4;
  input [20:5] PP5;
  input [21:6] PP6;
  input [22:7] PP7;
  input [23:8] PP8;
  input [24:9] PP9;
  wire [29:6] W0;
  wire [31:0] W1;
  wire [30:3] W2;
  OSBODY_15_0_16_1_000 U0 (W0, W1, W2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15);
  CSA_29_6_31_0_30_000 U1 (S1, S2, W0, W1, W2);
endmodule

module PureCSA_15_2 (C, S, X, Y, Z);
  output [16:3] C;
  output [15:2] S;
  input [15:2] X;
  input [15:2] Y;
  input [15:2] Z;
  UBFA_2 U0 (C[3], S[2], X[2], Y[2], Z[2]);
  UBFA_3 U1 (C[4], S[3], X[3], Y[3], Z[3]);
  UBFA_4 U2 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U3 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U4 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U5 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U6 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U7 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U8 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U9 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U10 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U11 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U12 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U13 (C[16], S[15], X[15], Y[15], Z[15]);
endmodule

module PureCSA_17_5 (C, S, X, Y, Z);
  output [18:6] C;
  output [17:5] S;
  input [17:5] X;
  input [17:5] Y;
  input [17:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U3 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U4 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U5 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U6 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U7 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U8 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U9 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U10 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U11 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U12 (C[18], S[17], X[17], Y[17], Z[17]);
endmodule

module PureCSA_18_5 (C, S, X, Y, Z);
  output [19:6] C;
  output [18:5] S;
  input [18:5] X;
  input [18:5] Y;
  input [18:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U3 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U4 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U5 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U6 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U7 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U8 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U9 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U10 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U11 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U12 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U13 (C[19], S[18], X[18], Y[18], Z[18]);
endmodule

module PureCSA_18_7 (C, S, X, Y, Z);
  output [19:8] C;
  output [18:7] S;
  input [18:7] X;
  input [18:7] Y;
  input [18:7] Z;
  UBFA_7 U0 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U1 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U2 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U3 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U4 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U5 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U6 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U7 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U8 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U9 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U10 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U11 (C[19], S[18], X[18], Y[18], Z[18]);
endmodule

module PureCSA_20_8 (C, S, X, Y, Z);
  output [21:9] C;
  output [20:8] S;
  input [20:8] X;
  input [20:8] Y;
  input [20:8] Z;
  UBFA_8 U0 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U1 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U2 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U3 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U4 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U5 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U6 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U7 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U8 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U9 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U10 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U11 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U12 (C[21], S[20], X[20], Y[20], Z[20]);
endmodule

module PureCSA_21_10 (C, S, X, Y, Z);
  output [22:11] C;
  output [21:10] S;
  input [21:10] X;
  input [21:10] Y;
  input [21:10] Z;
  UBFA_10 U0 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U1 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U2 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U3 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U4 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U5 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U6 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U7 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U8 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U9 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U10 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U11 (C[22], S[21], X[21], Y[21], Z[21]);
endmodule

module PureCSA_21_8 (C, S, X, Y, Z);
  output [22:9] C;
  output [21:8] S;
  input [21:8] X;
  input [21:8] Y;
  input [21:8] Z;
  UBFA_8 U0 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U1 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U2 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U3 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U4 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U5 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U6 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U7 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U8 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U9 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U10 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U11 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U12 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U13 (C[22], S[21], X[21], Y[21], Z[21]);
endmodule

module PureCSA_23_12 (C, S, X, Y, Z);
  output [24:13] C;
  output [23:12] S;
  input [23:12] X;
  input [23:12] Y;
  input [23:12] Z;
  UBFA_12 U0 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U1 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U2 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U3 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U4 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U5 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U6 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U7 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U8 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U9 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U10 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U11 (C[24], S[23], X[23], Y[23], Z[23]);
endmodule

module PureCSA_24_11 (C, S, X, Y, Z);
  output [25:12] C;
  output [24:11] S;
  input [24:11] X;
  input [24:11] Y;
  input [24:11] Z;
  UBFA_11 U0 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U1 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U2 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U3 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U4 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U5 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U6 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U7 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U8 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U9 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U10 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U11 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U12 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U13 (C[25], S[24], X[24], Y[24], Z[24]);
endmodule

module PureCSA_25_14 (C, S, X, Y, Z);
  output [26:15] C;
  output [25:14] S;
  input [25:14] X;
  input [25:14] Y;
  input [25:14] Z;
  UBFA_14 U0 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U1 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U2 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U3 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U4 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U5 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U6 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U7 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U8 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U9 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U10 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U11 (C[26], S[25], X[25], Y[25], Z[25]);
endmodule

module PureCSA_26_12 (C, S, X, Y, Z);
  output [27:13] C;
  output [26:12] S;
  input [26:12] X;
  input [26:12] Y;
  input [26:12] Z;
  UBFA_12 U0 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U1 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U2 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U3 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U4 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U5 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U6 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U7 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U8 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U9 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U10 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U11 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U12 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U13 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U14 (C[27], S[26], X[26], Y[26], Z[26]);
endmodule

module PureCSA_27_15 (C, S, X, Y, Z);
  output [28:16] C;
  output [27:15] S;
  input [27:15] X;
  input [27:15] Y;
  input [27:15] Z;
  UBFA_15 U0 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U1 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U2 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U3 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U4 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U5 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U6 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U7 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U8 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U9 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U10 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U11 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U12 (C[28], S[27], X[27], Y[27], Z[27]);
endmodule

module PureCSA_28_15 (C, S, X, Y, Z);
  output [29:16] C;
  output [28:15] S;
  input [28:15] X;
  input [28:15] Y;
  input [28:15] Z;
  UBFA_15 U0 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U1 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U2 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U3 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U4 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U5 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U6 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U7 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U8 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U9 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U10 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U11 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U12 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U13 (C[29], S[28], X[28], Y[28], Z[28]);
endmodule

module PureCSA_29_6 (C, S, X, Y, Z);
  output [30:7] C;
  output [29:6] S;
  input [29:6] X;
  input [29:6] Y;
  input [29:6] Z;
  UBFA_6 U0 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U1 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U2 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U3 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U4 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U5 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U6 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U7 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U8 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U9 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U10 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U11 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U12 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U13 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U14 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U15 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U16 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U17 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U18 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U19 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U20 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U21 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U22 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U23 (C[30], S[29], X[29], Y[29], Z[29]);
endmodule

module PureCSHA_11_9 (C, S, X, Y);
  output [12:10] C;
  output [11:9] S;
  input [11:9] X;
  input [11:9] Y;
  UBHA_9 U0 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U1 (C[11], S[10], X[10], Y[10]);
  UBHA_11 U2 (C[12], S[11], X[11], Y[11]);
endmodule

module PureCSHA_13_5 (C, S, X, Y);
  output [14:6] C;
  output [13:5] S;
  input [13:5] X;
  input [13:5] Y;
  UBHA_5 U0 (C[6], S[5], X[5], Y[5]);
  UBHA_6 U1 (C[7], S[6], X[6], Y[6]);
  UBHA_7 U2 (C[8], S[7], X[7], Y[7]);
  UBHA_8 U3 (C[9], S[8], X[8], Y[8]);
  UBHA_9 U4 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U5 (C[11], S[10], X[10], Y[10]);
  UBHA_11 U6 (C[12], S[11], X[11], Y[11]);
  UBHA_12 U7 (C[13], S[12], X[12], Y[12]);
  UBHA_13 U8 (C[14], S[13], X[13], Y[13]);
endmodule

module PureCSHA_14_13 (C, S, X, Y);
  output [15:14] C;
  output [14:13] S;
  input [14:13] X;
  input [14:13] Y;
  UBHA_13 U0 (C[14], S[13], X[13], Y[13]);
  UBHA_14 U1 (C[15], S[14], X[14], Y[14]);
endmodule

module PureCSHA_20_19 (C, S, X, Y);
  output [21:20] C;
  output [20:19] S;
  input [20:19] X;
  input [20:19] Y;
  UBHA_19 U0 (C[20], S[19], X[19], Y[19]);
  UBHA_20 U1 (C[21], S[20], X[20], Y[20]);
endmodule

module PureCSHA_23_21 (C, S, X, Y);
  output [24:22] C;
  output [23:21] S;
  input [23:21] X;
  input [23:21] Y;
  UBHA_21 U0 (C[22], S[21], X[21], Y[21]);
  UBHA_22 U1 (C[23], S[22], X[22], Y[22]);
  UBHA_23 U2 (C[24], S[23], X[23], Y[23]);
endmodule

module PureCSHA_24_22 (C, S, X, Y);
  output [25:23] C;
  output [24:22] S;
  input [24:22] X;
  input [24:22] Y;
  UBHA_22 U0 (C[23], S[22], X[22], Y[22]);
  UBHA_23 U1 (C[24], S[23], X[23], Y[23]);
  UBHA_24 U2 (C[25], S[24], X[24], Y[24]);
endmodule

module PureCSHA_27_24 (C, S, X, Y);
  output [28:25] C;
  output [27:24] S;
  input [27:24] X;
  input [27:24] Y;
  UBHA_24 U0 (C[25], S[24], X[24], Y[24]);
  UBHA_25 U1 (C[26], S[25], X[25], Y[25]);
  UBHA_26 U2 (C[27], S[26], X[26], Y[26]);
  UBHA_27 U3 (C[28], S[27], X[27], Y[27]);
endmodule

module PureCSHA_28_26 (C, S, X, Y);
  output [29:27] C;
  output [28:26] S;
  input [28:26] X;
  input [28:26] Y;
  UBHA_26 U0 (C[27], S[26], X[26], Y[26]);
  UBHA_27 U1 (C[28], S[27], X[27], Y[27]);
  UBHA_28 U2 (C[29], S[28], X[28], Y[28]);
endmodule

module PureCSHA_30_28 (C, S, X, Y);
  output [31:29] C;
  output [30:28] S;
  input [30:28] X;
  input [30:28] Y;
  UBHA_28 U0 (C[29], S[28], X[28], Y[28]);
  UBHA_29 U1 (C[30], S[29], X[29], Y[29]);
  UBHA_30 U2 (C[31], S[30], X[30], Y[30]);
endmodule

module PureCSHA_4_2 (C, S, X, Y);
  output [5:3] C;
  output [4:2] S;
  input [4:2] X;
  input [4:2] Y;
  UBHA_2 U0 (C[3], S[2], X[2], Y[2]);
  UBHA_3 U1 (C[4], S[3], X[3], Y[3]);
  UBHA_4 U2 (C[5], S[4], X[4], Y[4]);
endmodule

module PureCSHA_5_3 (C, S, X, Y);
  output [6:4] C;
  output [5:3] S;
  input [5:3] X;
  input [5:3] Y;
  UBHA_3 U0 (C[4], S[3], X[3], Y[3]);
  UBHA_4 U1 (C[5], S[4], X[4], Y[4]);
  UBHA_5 U2 (C[6], S[5], X[5], Y[5]);
endmodule

module PureCSHA_6_3 (C, S, X, Y);
  output [7:4] C;
  output [6:3] S;
  input [6:3] X;
  input [6:3] Y;
  UBHA_3 U0 (C[4], S[3], X[3], Y[3]);
  UBHA_4 U1 (C[5], S[4], X[4], Y[4]);
  UBHA_5 U2 (C[6], S[5], X[5], Y[5]);
  UBHA_6 U3 (C[7], S[6], X[6], Y[6]);
endmodule

module PureCSHA_7_6 (C, S, X, Y);
  output [8:7] C;
  output [7:6] S;
  input [7:6] X;
  input [7:6] Y;
  UBHA_6 U0 (C[7], S[6], X[6], Y[6]);
  UBHA_7 U1 (C[8], S[7], X[7], Y[7]);
endmodule

module PureCSHA_9_4 (C, S, X, Y);
  output [10:5] C;
  output [9:4] S;
  input [9:4] X;
  input [9:4] Y;
  UBHA_4 U0 (C[5], S[4], X[4], Y[4]);
  UBHA_5 U1 (C[6], S[5], X[5], Y[5]);
  UBHA_6 U2 (C[7], S[6], X[6], Y[6]);
  UBHA_7 U3 (C[8], S[7], X[7], Y[7]);
  UBHA_8 U4 (C[9], S[8], X[8], Y[8]);
  UBHA_9 U5 (C[10], S[9], X[9], Y[9]);
endmodule

module UBARYACC_19_4_20_000 (S1, S2, PP0, PP1);
  output [19:4] S1;
  output [20:5] S2;
  input [19:4] PP0;
  input [20:5] PP1;
  UBCON_19_4 U0 (S1, PP0);
  UBCON_20_5 U1 (S2, PP1);
endmodule

module UBARYACC_21_6_22_000 (S1, S2, PP0, PP1, PP2);
  output [23:8] S1;
  output [23:6] S2;
  input [21:6] PP0;
  input [22:7] PP1;
  input [23:8] PP2;
  CSA_21_6_22_7_23_000 U0 (S1, S2, PP0, PP1, PP2);
endmodule

module UBARYACC_24_9_25_000 (S1, S2, PP0, PP1, PP2, PP3);
  output [27:12] S1;
  output [27:9] S2;
  input [24:9] PP0;
  input [25:10] PP1;
  input [26:11] PP2;
  input [27:12] PP3;
  wire [26:11] IC0;
  wire [26:9] IS0;
  CSA_24_9_25_10_26000 U0 (IC0, IS0, PP0, PP1, PP2);
  CSA_26_9_26_11_27000 U1 (S1, S2, IS0, IC0, PP3);
endmodule

module UBARYACC_28_13_29000 (S1, S2, PP0, PP1, PP2);
  output [30:15] S1;
  output [30:13] S2;
  input [28:13] PP0;
  input [29:14] PP1;
  input [30:15] PP2;
  CSA_28_13_29_14_3000 U0 (S1, S2, PP0, PP1, PP2);
endmodule

module UBCON_10_9 (O, I);
  output [10:9] O;
  input [10:9] I;
  UB1DCON_9 U0 (O[9], I[9]);
  UB1DCON_10 U1 (O[10], I[10]);
endmodule

module UBCON_12_3 (O, I);
  output [12:3] O;
  input [12:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
  UB1DCON_6 U3 (O[6], I[6]);
  UB1DCON_7 U4 (O[7], I[7]);
  UB1DCON_8 U5 (O[8], I[8]);
  UB1DCON_9 U6 (O[9], I[9]);
  UB1DCON_10 U7 (O[10], I[10]);
  UB1DCON_11 U8 (O[11], I[11]);
  UB1DCON_12 U9 (O[12], I[12]);
endmodule

module UBCON_18_3 (O, I);
  output [18:3] O;
  input [18:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
  UB1DCON_6 U3 (O[6], I[6]);
  UB1DCON_7 U4 (O[7], I[7]);
  UB1DCON_8 U5 (O[8], I[8]);
  UB1DCON_9 U6 (O[9], I[9]);
  UB1DCON_10 U7 (O[10], I[10]);
  UB1DCON_11 U8 (O[11], I[11]);
  UB1DCON_12 U9 (O[12], I[12]);
  UB1DCON_13 U10 (O[13], I[13]);
  UB1DCON_14 U11 (O[14], I[14]);
  UB1DCON_15 U12 (O[15], I[15]);
  UB1DCON_16 U13 (O[16], I[16]);
  UB1DCON_17 U14 (O[17], I[17]);
  UB1DCON_18 U15 (O[18], I[18]);
endmodule

module UBCON_19_4 (O, I);
  output [19:4] O;
  input [19:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
  UB1DCON_11 U7 (O[11], I[11]);
  UB1DCON_12 U8 (O[12], I[12]);
  UB1DCON_13 U9 (O[13], I[13]);
  UB1DCON_14 U10 (O[14], I[14]);
  UB1DCON_15 U11 (O[15], I[15]);
  UB1DCON_16 U12 (O[16], I[16]);
  UB1DCON_17 U13 (O[17], I[17]);
  UB1DCON_18 U14 (O[18], I[18]);
  UB1DCON_19 U15 (O[19], I[19]);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_20_18 (O, I);
  output [20:18] O;
  input [20:18] I;
  UB1DCON_18 U0 (O[18], I[18]);
  UB1DCON_19 U1 (O[19], I[19]);
  UB1DCON_20 U2 (O[20], I[20]);
endmodule

module UBCON_20_5 (O, I);
  output [20:5] O;
  input [20:5] I;
  UB1DCON_5 U0 (O[5], I[5]);
  UB1DCON_6 U1 (O[6], I[6]);
  UB1DCON_7 U2 (O[7], I[7]);
  UB1DCON_8 U3 (O[8], I[8]);
  UB1DCON_9 U4 (O[9], I[9]);
  UB1DCON_10 U5 (O[10], I[10]);
  UB1DCON_11 U6 (O[11], I[11]);
  UB1DCON_12 U7 (O[12], I[12]);
  UB1DCON_13 U8 (O[13], I[13]);
  UB1DCON_14 U9 (O[14], I[14]);
  UB1DCON_15 U10 (O[15], I[15]);
  UB1DCON_16 U11 (O[16], I[16]);
  UB1DCON_17 U12 (O[17], I[17]);
  UB1DCON_18 U13 (O[18], I[18]);
  UB1DCON_19 U14 (O[19], I[19]);
  UB1DCON_20 U15 (O[20], I[20]);
endmodule

module UBCON_24_21 (O, I);
  output [24:21] O;
  input [24:21] I;
  UB1DCON_21 U0 (O[21], I[21]);
  UB1DCON_22 U1 (O[22], I[22]);
  UB1DCON_23 U2 (O[23], I[23]);
  UB1DCON_24 U3 (O[24], I[24]);
endmodule

module UBCON_28_25 (O, I);
  output [28:25] O;
  input [28:25] I;
  UB1DCON_25 U0 (O[25], I[25]);
  UB1DCON_26 U1 (O[26], I[26]);
  UB1DCON_27 U2 (O[27], I[27]);
  UB1DCON_28 U3 (O[28], I[28]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBCON_31_29 (O, I);
  output [31:29] O;
  input [31:29] I;
  UB1DCON_29 U0 (O[29], I[29]);
  UB1DCON_30 U1 (O[30], I[30]);
  UB1DCON_31 U2 (O[31], I[31]);
endmodule

module UBCON_3_0 (O, I);
  output [3:0] O;
  input [3:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
endmodule

module UBCON_4_0 (O, I);
  output [4:0] O;
  input [4:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
endmodule

module UBCON_5_3 (O, I);
  output [5:3] O;
  input [5:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
endmodule

module UBCON_8_3 (O, I);
  output [8:3] O;
  input [8:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
  UB1DCON_6 U3 (O[6], I[6]);
  UB1DCON_7 U4 (O[7], I[7]);
  UB1DCON_8 U5 (O[8], I[8]);
endmodule

module UBFCSkA_31_4_31_0 (S, X, Y);
  output [32:0] S;
  input [31:4] X;
  input [31:0] Y;
  UBPureFCSkA_31_4 U0 (S[32:4], X[31:4], Y[31:4]);
  UBCON_3_0 U1 (S[3:0], Y[3:0]);
endmodule

module UBPPG_15_0_15_0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, IN1, IN2);
  output [15:0] PP0;
  output [16:1] PP1;
  output [25:10] PP10;
  output [26:11] PP11;
  output [27:12] PP12;
  output [28:13] PP13;
  output [29:14] PP14;
  output [30:15] PP15;
  output [17:2] PP2;
  output [18:3] PP3;
  output [19:4] PP4;
  output [20:5] PP5;
  output [21:6] PP6;
  output [22:7] PP7;
  output [23:8] PP8;
  output [24:9] PP9;
  input [15:0] IN1;
  input [15:0] IN2;
  UBVPPG_15_0_0 U0 (PP0, IN1, IN2[0]);
  UBVPPG_15_0_1 U1 (PP1, IN1, IN2[1]);
  UBVPPG_15_0_2 U2 (PP2, IN1, IN2[2]);
  UBVPPG_15_0_3 U3 (PP3, IN1, IN2[3]);
  UBVPPG_15_0_4 U4 (PP4, IN1, IN2[4]);
  UBVPPG_15_0_5 U5 (PP5, IN1, IN2[5]);
  UBVPPG_15_0_6 U6 (PP6, IN1, IN2[6]);
  UBVPPG_15_0_7 U7 (PP7, IN1, IN2[7]);
  UBVPPG_15_0_8 U8 (PP8, IN1, IN2[8]);
  UBVPPG_15_0_9 U9 (PP9, IN1, IN2[9]);
  UBVPPG_15_0_10 U10 (PP10, IN1, IN2[10]);
  UBVPPG_15_0_11 U11 (PP11, IN1, IN2[11]);
  UBVPPG_15_0_12 U12 (PP12, IN1, IN2[12]);
  UBVPPG_15_0_13 U13 (PP13, IN1, IN2[13]);
  UBVPPG_15_0_14 U14 (PP14, IN1, IN2[14]);
  UBVPPG_15_0_15 U15 (PP15, IN1, IN2[15]);
endmodule

module UBPureFCSkA_31_4 (S, X, Y);
  output [32:4] S;
  input [31:4] X;
  input [31:4] Y;
  wire C;
  UBPriFCSkA_31_4 U0 (S, X, Y, C);
  UBZero_4_4 U1 (C);
endmodule

module UBVPPG_15_0_0 (O, IN1, IN2);
  output [15:0] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
  UB1BPPG_6_0 U6 (O[6], IN1[6], IN2);
  UB1BPPG_7_0 U7 (O[7], IN1[7], IN2);
  UB1BPPG_8_0 U8 (O[8], IN1[8], IN2);
  UB1BPPG_9_0 U9 (O[9], IN1[9], IN2);
  UB1BPPG_10_0 U10 (O[10], IN1[10], IN2);
  UB1BPPG_11_0 U11 (O[11], IN1[11], IN2);
  UB1BPPG_12_0 U12 (O[12], IN1[12], IN2);
  UB1BPPG_13_0 U13 (O[13], IN1[13], IN2);
  UB1BPPG_14_0 U14 (O[14], IN1[14], IN2);
  UB1BPPG_15_0 U15 (O[15], IN1[15], IN2);
endmodule

module UBVPPG_15_0_1 (O, IN1, IN2);
  output [16:1] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_1 U0 (O[1], IN1[0], IN2);
  UB1BPPG_1_1 U1 (O[2], IN1[1], IN2);
  UB1BPPG_2_1 U2 (O[3], IN1[2], IN2);
  UB1BPPG_3_1 U3 (O[4], IN1[3], IN2);
  UB1BPPG_4_1 U4 (O[5], IN1[4], IN2);
  UB1BPPG_5_1 U5 (O[6], IN1[5], IN2);
  UB1BPPG_6_1 U6 (O[7], IN1[6], IN2);
  UB1BPPG_7_1 U7 (O[8], IN1[7], IN2);
  UB1BPPG_8_1 U8 (O[9], IN1[8], IN2);
  UB1BPPG_9_1 U9 (O[10], IN1[9], IN2);
  UB1BPPG_10_1 U10 (O[11], IN1[10], IN2);
  UB1BPPG_11_1 U11 (O[12], IN1[11], IN2);
  UB1BPPG_12_1 U12 (O[13], IN1[12], IN2);
  UB1BPPG_13_1 U13 (O[14], IN1[13], IN2);
  UB1BPPG_14_1 U14 (O[15], IN1[14], IN2);
  UB1BPPG_15_1 U15 (O[16], IN1[15], IN2);
endmodule

module UBVPPG_15_0_10 (O, IN1, IN2);
  output [25:10] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_10 U0 (O[10], IN1[0], IN2);
  UB1BPPG_1_10 U1 (O[11], IN1[1], IN2);
  UB1BPPG_2_10 U2 (O[12], IN1[2], IN2);
  UB1BPPG_3_10 U3 (O[13], IN1[3], IN2);
  UB1BPPG_4_10 U4 (O[14], IN1[4], IN2);
  UB1BPPG_5_10 U5 (O[15], IN1[5], IN2);
  UB1BPPG_6_10 U6 (O[16], IN1[6], IN2);
  UB1BPPG_7_10 U7 (O[17], IN1[7], IN2);
  UB1BPPG_8_10 U8 (O[18], IN1[8], IN2);
  UB1BPPG_9_10 U9 (O[19], IN1[9], IN2);
  UB1BPPG_10_10 U10 (O[20], IN1[10], IN2);
  UB1BPPG_11_10 U11 (O[21], IN1[11], IN2);
  UB1BPPG_12_10 U12 (O[22], IN1[12], IN2);
  UB1BPPG_13_10 U13 (O[23], IN1[13], IN2);
  UB1BPPG_14_10 U14 (O[24], IN1[14], IN2);
  UB1BPPG_15_10 U15 (O[25], IN1[15], IN2);
endmodule

module UBVPPG_15_0_11 (O, IN1, IN2);
  output [26:11] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_11 U0 (O[11], IN1[0], IN2);
  UB1BPPG_1_11 U1 (O[12], IN1[1], IN2);
  UB1BPPG_2_11 U2 (O[13], IN1[2], IN2);
  UB1BPPG_3_11 U3 (O[14], IN1[3], IN2);
  UB1BPPG_4_11 U4 (O[15], IN1[4], IN2);
  UB1BPPG_5_11 U5 (O[16], IN1[5], IN2);
  UB1BPPG_6_11 U6 (O[17], IN1[6], IN2);
  UB1BPPG_7_11 U7 (O[18], IN1[7], IN2);
  UB1BPPG_8_11 U8 (O[19], IN1[8], IN2);
  UB1BPPG_9_11 U9 (O[20], IN1[9], IN2);
  UB1BPPG_10_11 U10 (O[21], IN1[10], IN2);
  UB1BPPG_11_11 U11 (O[22], IN1[11], IN2);
  UB1BPPG_12_11 U12 (O[23], IN1[12], IN2);
  UB1BPPG_13_11 U13 (O[24], IN1[13], IN2);
  UB1BPPG_14_11 U14 (O[25], IN1[14], IN2);
  UB1BPPG_15_11 U15 (O[26], IN1[15], IN2);
endmodule

module UBVPPG_15_0_12 (O, IN1, IN2);
  output [27:12] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_12 U0 (O[12], IN1[0], IN2);
  UB1BPPG_1_12 U1 (O[13], IN1[1], IN2);
  UB1BPPG_2_12 U2 (O[14], IN1[2], IN2);
  UB1BPPG_3_12 U3 (O[15], IN1[3], IN2);
  UB1BPPG_4_12 U4 (O[16], IN1[4], IN2);
  UB1BPPG_5_12 U5 (O[17], IN1[5], IN2);
  UB1BPPG_6_12 U6 (O[18], IN1[6], IN2);
  UB1BPPG_7_12 U7 (O[19], IN1[7], IN2);
  UB1BPPG_8_12 U8 (O[20], IN1[8], IN2);
  UB1BPPG_9_12 U9 (O[21], IN1[9], IN2);
  UB1BPPG_10_12 U10 (O[22], IN1[10], IN2);
  UB1BPPG_11_12 U11 (O[23], IN1[11], IN2);
  UB1BPPG_12_12 U12 (O[24], IN1[12], IN2);
  UB1BPPG_13_12 U13 (O[25], IN1[13], IN2);
  UB1BPPG_14_12 U14 (O[26], IN1[14], IN2);
  UB1BPPG_15_12 U15 (O[27], IN1[15], IN2);
endmodule

module UBVPPG_15_0_13 (O, IN1, IN2);
  output [28:13] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_13 U0 (O[13], IN1[0], IN2);
  UB1BPPG_1_13 U1 (O[14], IN1[1], IN2);
  UB1BPPG_2_13 U2 (O[15], IN1[2], IN2);
  UB1BPPG_3_13 U3 (O[16], IN1[3], IN2);
  UB1BPPG_4_13 U4 (O[17], IN1[4], IN2);
  UB1BPPG_5_13 U5 (O[18], IN1[5], IN2);
  UB1BPPG_6_13 U6 (O[19], IN1[6], IN2);
  UB1BPPG_7_13 U7 (O[20], IN1[7], IN2);
  UB1BPPG_8_13 U8 (O[21], IN1[8], IN2);
  UB1BPPG_9_13 U9 (O[22], IN1[9], IN2);
  UB1BPPG_10_13 U10 (O[23], IN1[10], IN2);
  UB1BPPG_11_13 U11 (O[24], IN1[11], IN2);
  UB1BPPG_12_13 U12 (O[25], IN1[12], IN2);
  UB1BPPG_13_13 U13 (O[26], IN1[13], IN2);
  UB1BPPG_14_13 U14 (O[27], IN1[14], IN2);
  UB1BPPG_15_13 U15 (O[28], IN1[15], IN2);
endmodule

module UBVPPG_15_0_14 (O, IN1, IN2);
  output [29:14] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_14 U0 (O[14], IN1[0], IN2);
  UB1BPPG_1_14 U1 (O[15], IN1[1], IN2);
  UB1BPPG_2_14 U2 (O[16], IN1[2], IN2);
  UB1BPPG_3_14 U3 (O[17], IN1[3], IN2);
  UB1BPPG_4_14 U4 (O[18], IN1[4], IN2);
  UB1BPPG_5_14 U5 (O[19], IN1[5], IN2);
  UB1BPPG_6_14 U6 (O[20], IN1[6], IN2);
  UB1BPPG_7_14 U7 (O[21], IN1[7], IN2);
  UB1BPPG_8_14 U8 (O[22], IN1[8], IN2);
  UB1BPPG_9_14 U9 (O[23], IN1[9], IN2);
  UB1BPPG_10_14 U10 (O[24], IN1[10], IN2);
  UB1BPPG_11_14 U11 (O[25], IN1[11], IN2);
  UB1BPPG_12_14 U12 (O[26], IN1[12], IN2);
  UB1BPPG_13_14 U13 (O[27], IN1[13], IN2);
  UB1BPPG_14_14 U14 (O[28], IN1[14], IN2);
  UB1BPPG_15_14 U15 (O[29], IN1[15], IN2);
endmodule

module UBVPPG_15_0_15 (O, IN1, IN2);
  output [30:15] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_15 U0 (O[15], IN1[0], IN2);
  UB1BPPG_1_15 U1 (O[16], IN1[1], IN2);
  UB1BPPG_2_15 U2 (O[17], IN1[2], IN2);
  UB1BPPG_3_15 U3 (O[18], IN1[3], IN2);
  UB1BPPG_4_15 U4 (O[19], IN1[4], IN2);
  UB1BPPG_5_15 U5 (O[20], IN1[5], IN2);
  UB1BPPG_6_15 U6 (O[21], IN1[6], IN2);
  UB1BPPG_7_15 U7 (O[22], IN1[7], IN2);
  UB1BPPG_8_15 U8 (O[23], IN1[8], IN2);
  UB1BPPG_9_15 U9 (O[24], IN1[9], IN2);
  UB1BPPG_10_15 U10 (O[25], IN1[10], IN2);
  UB1BPPG_11_15 U11 (O[26], IN1[11], IN2);
  UB1BPPG_12_15 U12 (O[27], IN1[12], IN2);
  UB1BPPG_13_15 U13 (O[28], IN1[13], IN2);
  UB1BPPG_14_15 U14 (O[29], IN1[14], IN2);
  UB1BPPG_15_15 U15 (O[30], IN1[15], IN2);
endmodule

module UBVPPG_15_0_2 (O, IN1, IN2);
  output [17:2] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
  UB1BPPG_6_2 U6 (O[8], IN1[6], IN2);
  UB1BPPG_7_2 U7 (O[9], IN1[7], IN2);
  UB1BPPG_8_2 U8 (O[10], IN1[8], IN2);
  UB1BPPG_9_2 U9 (O[11], IN1[9], IN2);
  UB1BPPG_10_2 U10 (O[12], IN1[10], IN2);
  UB1BPPG_11_2 U11 (O[13], IN1[11], IN2);
  UB1BPPG_12_2 U12 (O[14], IN1[12], IN2);
  UB1BPPG_13_2 U13 (O[15], IN1[13], IN2);
  UB1BPPG_14_2 U14 (O[16], IN1[14], IN2);
  UB1BPPG_15_2 U15 (O[17], IN1[15], IN2);
endmodule

module UBVPPG_15_0_3 (O, IN1, IN2);
  output [18:3] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_3 U0 (O[3], IN1[0], IN2);
  UB1BPPG_1_3 U1 (O[4], IN1[1], IN2);
  UB1BPPG_2_3 U2 (O[5], IN1[2], IN2);
  UB1BPPG_3_3 U3 (O[6], IN1[3], IN2);
  UB1BPPG_4_3 U4 (O[7], IN1[4], IN2);
  UB1BPPG_5_3 U5 (O[8], IN1[5], IN2);
  UB1BPPG_6_3 U6 (O[9], IN1[6], IN2);
  UB1BPPG_7_3 U7 (O[10], IN1[7], IN2);
  UB1BPPG_8_3 U8 (O[11], IN1[8], IN2);
  UB1BPPG_9_3 U9 (O[12], IN1[9], IN2);
  UB1BPPG_10_3 U10 (O[13], IN1[10], IN2);
  UB1BPPG_11_3 U11 (O[14], IN1[11], IN2);
  UB1BPPG_12_3 U12 (O[15], IN1[12], IN2);
  UB1BPPG_13_3 U13 (O[16], IN1[13], IN2);
  UB1BPPG_14_3 U14 (O[17], IN1[14], IN2);
  UB1BPPG_15_3 U15 (O[18], IN1[15], IN2);
endmodule

module UBVPPG_15_0_4 (O, IN1, IN2);
  output [19:4] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
  UB1BPPG_6_4 U6 (O[10], IN1[6], IN2);
  UB1BPPG_7_4 U7 (O[11], IN1[7], IN2);
  UB1BPPG_8_4 U8 (O[12], IN1[8], IN2);
  UB1BPPG_9_4 U9 (O[13], IN1[9], IN2);
  UB1BPPG_10_4 U10 (O[14], IN1[10], IN2);
  UB1BPPG_11_4 U11 (O[15], IN1[11], IN2);
  UB1BPPG_12_4 U12 (O[16], IN1[12], IN2);
  UB1BPPG_13_4 U13 (O[17], IN1[13], IN2);
  UB1BPPG_14_4 U14 (O[18], IN1[14], IN2);
  UB1BPPG_15_4 U15 (O[19], IN1[15], IN2);
endmodule

module UBVPPG_15_0_5 (O, IN1, IN2);
  output [20:5] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_5 U0 (O[5], IN1[0], IN2);
  UB1BPPG_1_5 U1 (O[6], IN1[1], IN2);
  UB1BPPG_2_5 U2 (O[7], IN1[2], IN2);
  UB1BPPG_3_5 U3 (O[8], IN1[3], IN2);
  UB1BPPG_4_5 U4 (O[9], IN1[4], IN2);
  UB1BPPG_5_5 U5 (O[10], IN1[5], IN2);
  UB1BPPG_6_5 U6 (O[11], IN1[6], IN2);
  UB1BPPG_7_5 U7 (O[12], IN1[7], IN2);
  UB1BPPG_8_5 U8 (O[13], IN1[8], IN2);
  UB1BPPG_9_5 U9 (O[14], IN1[9], IN2);
  UB1BPPG_10_5 U10 (O[15], IN1[10], IN2);
  UB1BPPG_11_5 U11 (O[16], IN1[11], IN2);
  UB1BPPG_12_5 U12 (O[17], IN1[12], IN2);
  UB1BPPG_13_5 U13 (O[18], IN1[13], IN2);
  UB1BPPG_14_5 U14 (O[19], IN1[14], IN2);
  UB1BPPG_15_5 U15 (O[20], IN1[15], IN2);
endmodule

module UBVPPG_15_0_6 (O, IN1, IN2);
  output [21:6] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_6 U0 (O[6], IN1[0], IN2);
  UB1BPPG_1_6 U1 (O[7], IN1[1], IN2);
  UB1BPPG_2_6 U2 (O[8], IN1[2], IN2);
  UB1BPPG_3_6 U3 (O[9], IN1[3], IN2);
  UB1BPPG_4_6 U4 (O[10], IN1[4], IN2);
  UB1BPPG_5_6 U5 (O[11], IN1[5], IN2);
  UB1BPPG_6_6 U6 (O[12], IN1[6], IN2);
  UB1BPPG_7_6 U7 (O[13], IN1[7], IN2);
  UB1BPPG_8_6 U8 (O[14], IN1[8], IN2);
  UB1BPPG_9_6 U9 (O[15], IN1[9], IN2);
  UB1BPPG_10_6 U10 (O[16], IN1[10], IN2);
  UB1BPPG_11_6 U11 (O[17], IN1[11], IN2);
  UB1BPPG_12_6 U12 (O[18], IN1[12], IN2);
  UB1BPPG_13_6 U13 (O[19], IN1[13], IN2);
  UB1BPPG_14_6 U14 (O[20], IN1[14], IN2);
  UB1BPPG_15_6 U15 (O[21], IN1[15], IN2);
endmodule

module UBVPPG_15_0_7 (O, IN1, IN2);
  output [22:7] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_7 U0 (O[7], IN1[0], IN2);
  UB1BPPG_1_7 U1 (O[8], IN1[1], IN2);
  UB1BPPG_2_7 U2 (O[9], IN1[2], IN2);
  UB1BPPG_3_7 U3 (O[10], IN1[3], IN2);
  UB1BPPG_4_7 U4 (O[11], IN1[4], IN2);
  UB1BPPG_5_7 U5 (O[12], IN1[5], IN2);
  UB1BPPG_6_7 U6 (O[13], IN1[6], IN2);
  UB1BPPG_7_7 U7 (O[14], IN1[7], IN2);
  UB1BPPG_8_7 U8 (O[15], IN1[8], IN2);
  UB1BPPG_9_7 U9 (O[16], IN1[9], IN2);
  UB1BPPG_10_7 U10 (O[17], IN1[10], IN2);
  UB1BPPG_11_7 U11 (O[18], IN1[11], IN2);
  UB1BPPG_12_7 U12 (O[19], IN1[12], IN2);
  UB1BPPG_13_7 U13 (O[20], IN1[13], IN2);
  UB1BPPG_14_7 U14 (O[21], IN1[14], IN2);
  UB1BPPG_15_7 U15 (O[22], IN1[15], IN2);
endmodule

module UBVPPG_15_0_8 (O, IN1, IN2);
  output [23:8] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_8 U0 (O[8], IN1[0], IN2);
  UB1BPPG_1_8 U1 (O[9], IN1[1], IN2);
  UB1BPPG_2_8 U2 (O[10], IN1[2], IN2);
  UB1BPPG_3_8 U3 (O[11], IN1[3], IN2);
  UB1BPPG_4_8 U4 (O[12], IN1[4], IN2);
  UB1BPPG_5_8 U5 (O[13], IN1[5], IN2);
  UB1BPPG_6_8 U6 (O[14], IN1[6], IN2);
  UB1BPPG_7_8 U7 (O[15], IN1[7], IN2);
  UB1BPPG_8_8 U8 (O[16], IN1[8], IN2);
  UB1BPPG_9_8 U9 (O[17], IN1[9], IN2);
  UB1BPPG_10_8 U10 (O[18], IN1[10], IN2);
  UB1BPPG_11_8 U11 (O[19], IN1[11], IN2);
  UB1BPPG_12_8 U12 (O[20], IN1[12], IN2);
  UB1BPPG_13_8 U13 (O[21], IN1[13], IN2);
  UB1BPPG_14_8 U14 (O[22], IN1[14], IN2);
  UB1BPPG_15_8 U15 (O[23], IN1[15], IN2);
endmodule

module UBVPPG_15_0_9 (O, IN1, IN2);
  output [24:9] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_9 U0 (O[9], IN1[0], IN2);
  UB1BPPG_1_9 U1 (O[10], IN1[1], IN2);
  UB1BPPG_2_9 U2 (O[11], IN1[2], IN2);
  UB1BPPG_3_9 U3 (O[12], IN1[3], IN2);
  UB1BPPG_4_9 U4 (O[13], IN1[4], IN2);
  UB1BPPG_5_9 U5 (O[14], IN1[5], IN2);
  UB1BPPG_6_9 U6 (O[15], IN1[6], IN2);
  UB1BPPG_7_9 U7 (O[16], IN1[7], IN2);
  UB1BPPG_8_9 U8 (O[17], IN1[8], IN2);
  UB1BPPG_9_9 U9 (O[18], IN1[9], IN2);
  UB1BPPG_10_9 U10 (O[19], IN1[10], IN2);
  UB1BPPG_11_9 U11 (O[20], IN1[11], IN2);
  UB1BPPG_12_9 U12 (O[21], IN1[12], IN2);
  UB1BPPG_13_9 U13 (O[22], IN1[13], IN2);
  UB1BPPG_14_9 U14 (O[23], IN1[14], IN2);
  UB1BPPG_15_9 U15 (O[24], IN1[15], IN2);
endmodule

