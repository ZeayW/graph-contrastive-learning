/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: Multiplier_13_0_1000

  Number system: Unsigned binary
  Multiplicand length: 14
  Multiplier length: 14
  Partial product generation: Simple PPG
  Partial product accumulation: Dadda tree
  Final stage addition: Block carry look-ahead adder
----------------------------------------------------------------------------*/

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UBHA_13(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_14(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_21(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_23(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_24(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_25(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_9(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_10(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_11(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_12(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_12(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_13(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_14(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_15(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_16(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_17(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_18(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_6(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_7(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_8(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_19(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_20(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_21(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_5(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_22(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_23(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_24(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_25(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module GPGenerator(Go, Po, A, B);
  output Go;
  output Po;
  input A;
  input B;
  assign Go = A & B;
  assign Po = A ^ B;
endmodule

module BCLAU_4(Go, Po, G, P, Cin);
  output Go;
  output Po;
  input Cin;
  input [3:0] G;
  input [3:0] P;
  assign Po = P[0] & P[1] & P[2] & P[3];
  assign Go = G[3] | ( P[3] & G[2] ) | ( P[3] & P[2] & G[1] ) | ( P[3] & P[2] & P[1] & G[0] );
endmodule

module BCLAlU_4(Go, Po, S, X, Y, Cin);
  output Go;
  output Po;
  output [3:0] S;
  input Cin;
  input [3:0] X;
  input [3:0] Y;
  wire [3:1] C;
  wire [3:0] G;
  wire [3:0] P;
  assign C[1] = G[0] | ( P[0] & Cin );
  assign C[2] = G[1] | ( P[1] & C[1] );
  assign C[3] = G[2] | ( P[2] & C[2] );
  assign S[0] = P[0] ^ Cin;
  assign S[1] = P[1] ^ C[1];
  assign S[2] = P[2] ^ C[2];
  assign S[3] = P[3] ^ C[3];
  GPGenerator U0 (G[0], P[0], X[0], Y[0]);
  GPGenerator U1 (G[1], P[1], X[1], Y[1]);
  GPGenerator U2 (G[2], P[2], X[2], Y[2]);
  GPGenerator U3 (G[3], P[3], X[3], Y[3]);
  BCLAU_4 U4 (Go, Po, G, P, Cin);
endmodule

module BCLAU_2(Go, Po, G, P, Cin);
  output Go;
  output Po;
  input Cin;
  input [1:0] G;
  input [1:0] P;
  assign Po = P[0] & P[1];
  assign Go = G[1] | ( P[1] & G[0] );
endmodule

module BCLAlU_2(Go, Po, S, X, Y, Cin);
  output Go;
  output Po;
  output [1:0] S;
  input Cin;
  input [1:0] X;
  input [1:0] Y;
  wire [1:1] C;
  wire [1:0] G;
  wire [1:0] P;
  assign C[1] = G[0] | ( P[0] & Cin );
  assign S[0] = P[0] ^ Cin;
  assign S[1] = P[1] ^ C[1];
  GPGenerator U0 (G[0], P[0], X[0], Y[0]);
  GPGenerator U1 (G[1], P[1], X[1], Y[1]);
  BCLAU_2 U2 (Go, Po, G, P, Cin);
endmodule

module BCLAU_3(Go, Po, G, P, Cin);
  output Go;
  output Po;
  input Cin;
  input [2:0] G;
  input [2:0] P;
  assign Po = P[0] & P[1] & P[2];
  assign Go = G[2] | ( P[2] & G[1] ) | ( P[2] & P[1] & G[0] );
endmodule

module PriMBCLA_26_1(S, X, Y, Cin);
  output [27:1] S;
  input Cin;
  input [26:1] X;
  input [26:1] Y;
  wire [6:0] C1;
  wire [1:0] C2;
  wire [6:0] G1;
  wire [1:0] G2;
  wire [6:0] P1;
  wire [1:0] P2;
  assign C1[0] = C2[0];
  assign C1[1] = G1[0] | ( P1[0] & C1[0] );
  assign C1[2] = G1[1] | ( P1[1] & C1[1] );
  assign C1[3] = G1[2] | ( P1[2] & C1[2] );
  assign C1[4] = C2[1];
  assign C1[5] = G1[4] | ( P1[4] & C1[4] );
  assign C1[6] = G1[5] | ( P1[5] & C1[5] );
  assign C2[0] = Cin;
  assign C2[1] = G2[0] | ( P2[0] & C2[0] );
  assign S[27] = G2[1] | ( P2[1] & C2[1] );
  BCLAlU_4 U0 (G1[0], P1[0], S[4:1], X[4:1], Y[4:1], C1[0]);
  BCLAlU_4 U1 (G1[1], P1[1], S[8:5], X[8:5], Y[8:5], C1[1]);
  BCLAlU_4 U2 (G1[2], P1[2], S[12:9], X[12:9], Y[12:9], C1[2]);
  BCLAlU_4 U3 (G1[3], P1[3], S[16:13], X[16:13], Y[16:13], C1[3]);
  BCLAlU_4 U4 (G1[4], P1[4], S[20:17], X[20:17], Y[20:17], C1[4]);
  BCLAlU_4 U5 (G1[5], P1[5], S[24:21], X[24:21], Y[24:21], C1[5]);
  BCLAlU_2 U6 (G1[6], P1[6], S[26:25], X[26:25], Y[26:25], C1[6]);
  BCLAU_4 U7 (G2[0], P2[0], G1[3:0], P1[3:0], C2[0]);
  BCLAU_3 U8 (G2[1], P2[1], G1[6:4], P1[6:4], C2[1]);
endmodule

module UBZero_1_1(O);
  output [1:1] O;
  assign O[1] = 0;
endmodule

module Multiplier_13_0_1000(P, IN1, IN2);
  output [27:0] P;
  input [13:0] IN1;
  input [13:0] IN2;
  wire [27:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  assign P[12] = W[12];
  assign P[13] = W[13];
  assign P[14] = W[14];
  assign P[15] = W[15];
  assign P[16] = W[16];
  assign P[17] = W[17];
  assign P[18] = W[18];
  assign P[19] = W[19];
  assign P[20] = W[20];
  assign P[21] = W[21];
  assign P[22] = W[22];
  assign P[23] = W[23];
  assign P[24] = W[24];
  assign P[25] = W[25];
  assign P[26] = W[26];
  assign P[27] = W[27];
  MultUB_STD_DAD_BC000 U0 (W, IN1, IN2);
endmodule

module DADTR_13_0_14_1_1000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13);
  output [26:0] S1;
  output [26:1] S2;
  input [13:0] PP0;
  input [14:1] PP1;
  input [23:10] PP10;
  input [24:11] PP11;
  input [25:12] PP12;
  input [26:13] PP13;
  input [15:2] PP2;
  input [16:3] PP3;
  input [17:4] PP4;
  input [18:5] PP5;
  input [19:6] PP6;
  input [20:7] PP7;
  input [21:8] PP8;
  input [22:9] PP9;
  wire [26:0] W0;
  wire [25:1] W1;
  wire [16:10] W10;
  wire [15:11] W11;
  wire [15:12] W12;
  wire [24:2] W2;
  wire [23:3] W3;
  wire [22:4] W4;
  wire [21:5] W5;
  wire [20:6] W6;
  wire [19:7] W7;
  wire [18:8] W8;
  wire [17:9] W9;
  UBHA_13 U0 (W11[14], W12[13], PP0[13], PP1[13]);
  UBHA_14 U1 (W12[15], W12[14], PP1[14], PP2[14]);
  UBCON_12_0 U2 (W0[12:0], PP0[12:0]);
  UB1DCON_13 U3 (W0[13], PP2[13]);
  UB1DCON_14 U4 (W0[14], PP3[14]);
  UB1DCON_15 U5 (W0[15], PP2[15]);
  UB1DCON_16 U6 (W0[16], PP3[16]);
  UB1DCON_17 U7 (W0[17], PP4[17]);
  UB1DCON_18 U8 (W0[18], PP5[18]);
  UB1DCON_19 U9 (W0[19], PP6[19]);
  UB1DCON_20 U10 (W0[20], PP7[20]);
  UB1DCON_21 U11 (W0[21], PP8[21]);
  UB1DCON_22 U12 (W0[22], PP9[22]);
  UB1DCON_23 U13 (W0[23], PP10[23]);
  UB1DCON_24 U14 (W0[24], PP11[24]);
  UB1DCON_25 U15 (W0[25], PP12[25]);
  UB1DCON_26 U16 (W0[26], PP13[26]);
  UBCON_12_1 U17 (W1[12:1], PP1[12:1]);
  UB1DCON_13 U18 (W1[13], PP3[13]);
  UB1DCON_14 U19 (W1[14], PP4[14]);
  UB1DCON_15 U20 (W1[15], PP3[15]);
  UB1DCON_16 U21 (W1[16], PP4[16]);
  UB1DCON_17 U22 (W1[17], PP5[17]);
  UB1DCON_18 U23 (W1[18], PP6[18]);
  UB1DCON_19 U24 (W1[19], PP7[19]);
  UB1DCON_20 U25 (W1[20], PP8[20]);
  UB1DCON_21 U26 (W1[21], PP9[21]);
  UB1DCON_22 U27 (W1[22], PP10[22]);
  UB1DCON_23 U28 (W1[23], PP11[23]);
  UB1DCON_24 U29 (W1[24], PP12[24]);
  UB1DCON_25 U30 (W1[25], PP13[25]);
  UBCON_12_2 U31 (W2[12:2], PP2[12:2]);
  UB1DCON_13 U32 (W2[13], PP4[13]);
  UB1DCON_14 U33 (W2[14], PP5[14]);
  UB1DCON_15 U34 (W2[15], PP4[15]);
  UB1DCON_16 U35 (W2[16], PP5[16]);
  UB1DCON_17 U36 (W2[17], PP6[17]);
  UB1DCON_18 U37 (W2[18], PP7[18]);
  UB1DCON_19 U38 (W2[19], PP8[19]);
  UB1DCON_20 U39 (W2[20], PP9[20]);
  UB1DCON_21 U40 (W2[21], PP10[21]);
  UB1DCON_22 U41 (W2[22], PP11[22]);
  UB1DCON_23 U42 (W2[23], PP12[23]);
  UB1DCON_24 U43 (W2[24], PP13[24]);
  UBCON_12_3 U44 (W3[12:3], PP3[12:3]);
  UB1DCON_13 U45 (W3[13], PP5[13]);
  UB1DCON_14 U46 (W3[14], PP6[14]);
  UB1DCON_15 U47 (W3[15], PP5[15]);
  UB1DCON_16 U48 (W3[16], PP6[16]);
  UB1DCON_17 U49 (W3[17], PP7[17]);
  UB1DCON_18 U50 (W3[18], PP8[18]);
  UB1DCON_19 U51 (W3[19], PP9[19]);
  UB1DCON_20 U52 (W3[20], PP10[20]);
  UB1DCON_21 U53 (W3[21], PP11[21]);
  UB1DCON_22 U54 (W3[22], PP12[22]);
  UB1DCON_23 U55 (W3[23], PP13[23]);
  UBCON_12_4 U56 (W4[12:4], PP4[12:4]);
  UB1DCON_13 U57 (W4[13], PP6[13]);
  UB1DCON_14 U58 (W4[14], PP7[14]);
  UB1DCON_15 U59 (W4[15], PP6[15]);
  UB1DCON_16 U60 (W4[16], PP7[16]);
  UB1DCON_17 U61 (W4[17], PP8[17]);
  UB1DCON_18 U62 (W4[18], PP9[18]);
  UB1DCON_19 U63 (W4[19], PP10[19]);
  UB1DCON_20 U64 (W4[20], PP11[20]);
  UB1DCON_21 U65 (W4[21], PP12[21]);
  UB1DCON_22 U66 (W4[22], PP13[22]);
  UBCON_12_5 U67 (W5[12:5], PP5[12:5]);
  UB1DCON_13 U68 (W5[13], PP7[13]);
  UB1DCON_14 U69 (W5[14], PP8[14]);
  UB1DCON_15 U70 (W5[15], PP7[15]);
  UB1DCON_16 U71 (W5[16], PP8[16]);
  UB1DCON_17 U72 (W5[17], PP9[17]);
  UB1DCON_18 U73 (W5[18], PP10[18]);
  UB1DCON_19 U74 (W5[19], PP11[19]);
  UB1DCON_20 U75 (W5[20], PP12[20]);
  UB1DCON_21 U76 (W5[21], PP13[21]);
  UBCON_12_6 U77 (W6[12:6], PP6[12:6]);
  UB1DCON_13 U78 (W6[13], PP8[13]);
  UB1DCON_14 U79 (W6[14], PP9[14]);
  UB1DCON_15 U80 (W6[15], PP8[15]);
  UB1DCON_16 U81 (W6[16], PP9[16]);
  UB1DCON_17 U82 (W6[17], PP10[17]);
  UB1DCON_18 U83 (W6[18], PP11[18]);
  UB1DCON_19 U84 (W6[19], PP12[19]);
  UB1DCON_20 U85 (W6[20], PP13[20]);
  UBCON_12_7 U86 (W7[12:7], PP7[12:7]);
  UB1DCON_13 U87 (W7[13], PP9[13]);
  UB1DCON_14 U88 (W7[14], PP10[14]);
  UB1DCON_15 U89 (W7[15], PP9[15]);
  UB1DCON_16 U90 (W7[16], PP10[16]);
  UB1DCON_17 U91 (W7[17], PP11[17]);
  UB1DCON_18 U92 (W7[18], PP12[18]);
  UB1DCON_19 U93 (W7[19], PP13[19]);
  UBCON_12_8 U94 (W8[12:8], PP8[12:8]);
  UB1DCON_13 U95 (W8[13], PP10[13]);
  UB1DCON_14 U96 (W8[14], PP11[14]);
  UB1DCON_15 U97 (W8[15], PP10[15]);
  UB1DCON_16 U98 (W8[16], PP11[16]);
  UB1DCON_17 U99 (W8[17], PP12[17]);
  UB1DCON_18 U100 (W8[18], PP13[18]);
  UBCON_12_9 U101 (W9[12:9], PP9[12:9]);
  UB1DCON_13 U102 (W9[13], PP11[13]);
  UB1DCON_14 U103 (W9[14], PP12[14]);
  UB1DCON_15 U104 (W9[15], PP11[15]);
  UB1DCON_16 U105 (W9[16], PP12[16]);
  UB1DCON_17 U106 (W9[17], PP13[17]);
  UBCON_12_10 U107 (W10[12:10], PP10[12:10]);
  UB1DCON_13 U108 (W10[13], PP12[13]);
  UB1DCON_14 U109 (W10[14], PP13[14]);
  UB1DCON_15 U110 (W10[15], PP12[15]);
  UB1DCON_16 U111 (W10[16], PP13[16]);
  UBCON_12_11 U112 (W11[12:11], PP11[12:11]);
  UB1DCON_13 U113 (W11[13], PP13[13]);
  UB1DCON_15 U114 (W11[15], PP13[15]);
  UB1DCON_12 U115 (W12[12], PP12[12]);
  DADTR_26_0_25_1_2000 U116 (S1, S2, W0, W1, W2, W3, W4, W5, W6, W7, W8, W9, W10, W11, W12);
endmodule

module DADTR_26_0_25_1_2000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12);
  output [26:0] S1;
  output [26:1] S2;
  input [26:0] PP0;
  input [25:1] PP1;
  input [16:10] PP10;
  input [15:11] PP11;
  input [15:12] PP12;
  input [24:2] PP2;
  input [23:3] PP3;
  input [22:4] PP4;
  input [21:5] PP5;
  input [20:6] PP6;
  input [19:7] PP7;
  input [18:8] PP8;
  input [17:9] PP9;
  wire [26:0] W0;
  wire [25:1] W1;
  wire [24:2] W2;
  wire [23:3] W3;
  wire [22:4] W4;
  wire [21:5] W5;
  wire [20:6] W6;
  wire [19:7] W7;
  wire [19:8] W8;
  UBHA_9 U0 (W6[10], W8[9], PP0[9], PP1[9]);
  UBFA_10 U1 (W4[11], W7[10], PP0[10], PP1[10], PP2[10]);
  UBHA_10 U2 (W5[11], W8[10], PP3[10], PP4[10]);
  UBFA_11 U3 (W2[12], W6[11], PP0[11], PP1[11], PP2[11]);
  UBFA_11 U4 (W3[12], W7[11], PP3[11], PP4[11], PP5[11]);
  UBHA_11 U5 (W4[12], W8[11], PP6[11], PP7[11]);
  UBFA_12 U6 (W1[13], W5[12], PP0[12], PP1[12], PP2[12]);
  UBFA_12 U7 (W2[13], W6[12], PP3[12], PP4[12], PP5[12]);
  UBFA_12 U8 (W3[13], W7[12], PP6[12], PP7[12], PP8[12]);
  UBHA_12 U9 (W4[13], W8[12], PP9[12], PP10[12]);
  UBFA_13 U10 (W1[14], W5[13], PP0[13], PP1[13], PP2[13]);
  UBFA_13 U11 (W2[14], W6[13], PP3[13], PP4[13], PP5[13]);
  UBFA_13 U12 (W3[14], W7[13], PP6[13], PP7[13], PP8[13]);
  UBFA_13 U13 (W4[14], W8[13], PP9[13], PP10[13], PP11[13]);
  UBFA_14 U14 (W1[15], W5[14], PP0[14], PP1[14], PP2[14]);
  UBFA_14 U15 (W2[15], W6[14], PP3[14], PP4[14], PP5[14]);
  UBFA_14 U16 (W3[15], W7[14], PP6[14], PP7[14], PP8[14]);
  UBFA_14 U17 (W4[15], W8[14], PP9[14], PP10[14], PP11[14]);
  UBFA_15 U18 (W2[16], W5[15], PP0[15], PP1[15], PP2[15]);
  UBFA_15 U19 (W3[16], W6[15], PP3[15], PP4[15], PP5[15]);
  UBFA_15 U20 (W4[16], W7[15], PP6[15], PP7[15], PP8[15]);
  UBFA_15 U21 (W5[16], W8[15], PP9[15], PP10[15], PP11[15]);
  UBFA_16 U22 (W4[17], W6[16], PP0[16], PP1[16], PP2[16]);
  UBFA_16 U23 (W5[17], W7[16], PP3[16], PP4[16], PP5[16]);
  UBFA_16 U24 (W6[17], W8[16], PP6[16], PP7[16], PP8[16]);
  UBFA_17 U25 (W6[18], W7[17], PP0[17], PP1[17], PP2[17]);
  UBFA_17 U26 (W7[18], W8[17], PP3[17], PP4[17], PP5[17]);
  UBFA_18 U27 (W8[19], W8[18], PP0[18], PP1[18], PP2[18]);
  UBCON_8_0 U28 (W0[8:0], PP0[8:0]);
  UB1DCON_9 U29 (W0[9], PP2[9]);
  UB1DCON_10 U30 (W0[10], PP5[10]);
  UB1DCON_11 U31 (W0[11], PP8[11]);
  UB1DCON_12 U32 (W0[12], PP11[12]);
  UBCON_15_13 U33 (W0[15:13], PP12[15:13]);
  UB1DCON_16 U34 (W0[16], PP9[16]);
  UB1DCON_17 U35 (W0[17], PP6[17]);
  UB1DCON_18 U36 (W0[18], PP3[18]);
  UBCON_26_19 U37 (W0[26:19], PP0[26:19]);
  UBCON_8_1 U38 (W1[8:1], PP1[8:1]);
  UB1DCON_9 U39 (W1[9], PP3[9]);
  UB1DCON_10 U40 (W1[10], PP6[10]);
  UB1DCON_11 U41 (W1[11], PP9[11]);
  UB1DCON_12 U42 (W1[12], PP12[12]);
  UB1DCON_16 U43 (W1[16], PP10[16]);
  UB1DCON_17 U44 (W1[17], PP7[17]);
  UB1DCON_18 U45 (W1[18], PP4[18]);
  UBCON_25_19 U46 (W1[25:19], PP1[25:19]);
  UBCON_8_2 U47 (W2[8:2], PP2[8:2]);
  UB1DCON_9 U48 (W2[9], PP4[9]);
  UB1DCON_10 U49 (W2[10], PP7[10]);
  UB1DCON_11 U50 (W2[11], PP10[11]);
  UB1DCON_17 U51 (W2[17], PP8[17]);
  UB1DCON_18 U52 (W2[18], PP5[18]);
  UBCON_24_19 U53 (W2[24:19], PP2[24:19]);
  UBCON_8_3 U54 (W3[8:3], PP3[8:3]);
  UB1DCON_9 U55 (W3[9], PP5[9]);
  UB1DCON_10 U56 (W3[10], PP8[10]);
  UB1DCON_11 U57 (W3[11], PP11[11]);
  UB1DCON_17 U58 (W3[17], PP9[17]);
  UB1DCON_18 U59 (W3[18], PP6[18]);
  UBCON_23_19 U60 (W3[23:19], PP3[23:19]);
  UBCON_8_4 U61 (W4[8:4], PP4[8:4]);
  UB1DCON_9 U62 (W4[9], PP6[9]);
  UB1DCON_10 U63 (W4[10], PP9[10]);
  UB1DCON_18 U64 (W4[18], PP7[18]);
  UBCON_22_19 U65 (W4[22:19], PP4[22:19]);
  UBCON_8_5 U66 (W5[8:5], PP5[8:5]);
  UB1DCON_9 U67 (W5[9], PP7[9]);
  UB1DCON_10 U68 (W5[10], PP10[10]);
  UB1DCON_18 U69 (W5[18], PP8[18]);
  UBCON_21_19 U70 (W5[21:19], PP5[21:19]);
  UBCON_8_6 U71 (W6[8:6], PP6[8:6]);
  UB1DCON_9 U72 (W6[9], PP8[9]);
  UBCON_20_19 U73 (W6[20:19], PP6[20:19]);
  UBCON_8_7 U74 (W7[8:7], PP7[8:7]);
  UB1DCON_9 U75 (W7[9], PP9[9]);
  UB1DCON_19 U76 (W7[19], PP7[19]);
  UB1DCON_8 U77 (W8[8], PP8[8]);
  DADTR_26_0_25_1_2001 U78 (S1, S2, W0, W1, W2, W3, W4, W5, W6, W7, W8);
endmodule

module DADTR_26_0_25_1_2001 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8);
  output [26:0] S1;
  output [26:1] S2;
  input [26:0] PP0;
  input [25:1] PP1;
  input [24:2] PP2;
  input [23:3] PP3;
  input [22:4] PP4;
  input [21:5] PP5;
  input [20:6] PP6;
  input [19:7] PP7;
  input [19:8] PP8;
  wire [26:0] W0;
  wire [25:1] W1;
  wire [24:2] W2;
  wire [23:3] W3;
  wire [22:4] W4;
  wire [22:5] W5;
  UBHA_6 U0 (W3[7], W5[6], PP0[6], PP1[6]);
  UBFA_7 U1 (W1[8], W4[7], PP0[7], PP1[7], PP2[7]);
  UBHA_7 U2 (W2[8], W5[7], PP3[7], PP4[7]);
  UBFA_8 U3 (W0[9], W3[8], PP0[8], PP1[8], PP2[8]);
  UBFA_8 U4 (W1[9], W4[8], PP3[8], PP4[8], PP5[8]);
  UBHA_8 U5 (W2[9], W5[8], PP6[8], PP7[8]);
  UBFA_9 U6 (W0[10], W3[9], PP0[9], PP1[9], PP2[9]);
  UBFA_9 U7 (W1[10], W4[9], PP3[9], PP4[9], PP5[9]);
  UBFA_9 U8 (W2[10], W5[9], PP6[9], PP7[9], PP8[9]);
  UBFA_10 U9 (W0[11], W3[10], PP0[10], PP1[10], PP2[10]);
  UBFA_10 U10 (W1[11], W4[10], PP3[10], PP4[10], PP5[10]);
  UBFA_10 U11 (W2[11], W5[10], PP6[10], PP7[10], PP8[10]);
  UBFA_11 U12 (W0[12], W3[11], PP0[11], PP1[11], PP2[11]);
  UBFA_11 U13 (W1[12], W4[11], PP3[11], PP4[11], PP5[11]);
  UBFA_11 U14 (W2[12], W5[11], PP6[11], PP7[11], PP8[11]);
  UBFA_12 U15 (W0[13], W3[12], PP0[12], PP1[12], PP2[12]);
  UBFA_12 U16 (W1[13], W4[12], PP3[12], PP4[12], PP5[12]);
  UBFA_12 U17 (W2[13], W5[12], PP6[12], PP7[12], PP8[12]);
  UBFA_13 U18 (W0[14], W3[13], PP0[13], PP1[13], PP2[13]);
  UBFA_13 U19 (W1[14], W4[13], PP3[13], PP4[13], PP5[13]);
  UBFA_13 U20 (W2[14], W5[13], PP6[13], PP7[13], PP8[13]);
  UBFA_14 U21 (W0[15], W3[14], PP0[14], PP1[14], PP2[14]);
  UBFA_14 U22 (W1[15], W4[14], PP3[14], PP4[14], PP5[14]);
  UBFA_14 U23 (W2[15], W5[14], PP6[14], PP7[14], PP8[14]);
  UBFA_15 U24 (W0[16], W3[15], PP0[15], PP1[15], PP2[15]);
  UBFA_15 U25 (W1[16], W4[15], PP3[15], PP4[15], PP5[15]);
  UBFA_15 U26 (W2[16], W5[15], PP6[15], PP7[15], PP8[15]);
  UBFA_16 U27 (W0[17], W3[16], PP0[16], PP1[16], PP2[16]);
  UBFA_16 U28 (W1[17], W4[16], PP3[16], PP4[16], PP5[16]);
  UBFA_16 U29 (W2[17], W5[16], PP6[16], PP7[16], PP8[16]);
  UBFA_17 U30 (W0[18], W3[17], PP0[17], PP1[17], PP2[17]);
  UBFA_17 U31 (W1[18], W4[17], PP3[17], PP4[17], PP5[17]);
  UBFA_17 U32 (W2[18], W5[17], PP6[17], PP7[17], PP8[17]);
  UBFA_18 U33 (W0[19], W3[18], PP0[18], PP1[18], PP2[18]);
  UBFA_18 U34 (W1[19], W4[18], PP3[18], PP4[18], PP5[18]);
  UBFA_18 U35 (W2[19], W5[18], PP6[18], PP7[18], PP8[18]);
  UBFA_19 U36 (W1[20], W3[19], PP0[19], PP1[19], PP2[19]);
  UBFA_19 U37 (W2[20], W4[19], PP3[19], PP4[19], PP5[19]);
  UBFA_19 U38 (W3[20], W5[19], PP6[19], PP7[19], PP8[19]);
  UBFA_20 U39 (W3[21], W4[20], PP0[20], PP1[20], PP2[20]);
  UBFA_20 U40 (W4[21], W5[20], PP3[20], PP4[20], PP5[20]);
  UBFA_21 U41 (W5[22], W5[21], PP0[21], PP1[21], PP2[21]);
  UBCON_5_0 U42 (W0[5:0], PP0[5:0]);
  UB1DCON_6 U43 (W0[6], PP2[6]);
  UB1DCON_7 U44 (W0[7], PP5[7]);
  UB1DCON_8 U45 (W0[8], PP8[8]);
  UB1DCON_20 U46 (W0[20], PP6[20]);
  UB1DCON_21 U47 (W0[21], PP3[21]);
  UBCON_26_22 U48 (W0[26:22], PP0[26:22]);
  UBCON_5_1 U49 (W1[5:1], PP1[5:1]);
  UB1DCON_6 U50 (W1[6], PP3[6]);
  UB1DCON_7 U51 (W1[7], PP6[7]);
  UB1DCON_21 U52 (W1[21], PP4[21]);
  UBCON_25_22 U53 (W1[25:22], PP1[25:22]);
  UBCON_5_2 U54 (W2[5:2], PP2[5:2]);
  UB1DCON_6 U55 (W2[6], PP4[6]);
  UB1DCON_7 U56 (W2[7], PP7[7]);
  UB1DCON_21 U57 (W2[21], PP5[21]);
  UBCON_24_22 U58 (W2[24:22], PP2[24:22]);
  UBCON_5_3 U59 (W3[5:3], PP3[5:3]);
  UB1DCON_6 U60 (W3[6], PP5[6]);
  UBCON_23_22 U61 (W3[23:22], PP3[23:22]);
  UBCON_5_4 U62 (W4[5:4], PP4[5:4]);
  UB1DCON_6 U63 (W4[6], PP6[6]);
  UB1DCON_22 U64 (W4[22], PP4[22]);
  UB1DCON_5 U65 (W5[5], PP5[5]);
  DADTR_26_0_25_1_2002 U66 (S1, S2, W0, W1, W2, W3, W4, W5);
endmodule

module DADTR_26_0_25_1_2002 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5);
  output [26:0] S1;
  output [26:1] S2;
  input [26:0] PP0;
  input [25:1] PP1;
  input [24:2] PP2;
  input [23:3] PP3;
  input [22:4] PP4;
  input [22:5] PP5;
  wire [26:0] W0;
  wire [25:1] W1;
  wire [24:2] W2;
  wire [24:3] W3;
  UBHA_4 U0 (W1[5], W3[4], PP0[4], PP1[4]);
  UBFA_5 U1 (W0[6], W2[5], PP0[5], PP1[5], PP2[5]);
  UBHA_5 U2 (W1[6], W3[5], PP3[5], PP4[5]);
  UBFA_6 U3 (W0[7], W2[6], PP0[6], PP1[6], PP2[6]);
  UBFA_6 U4 (W1[7], W3[6], PP3[6], PP4[6], PP5[6]);
  UBFA_7 U5 (W0[8], W2[7], PP0[7], PP1[7], PP2[7]);
  UBFA_7 U6 (W1[8], W3[7], PP3[7], PP4[7], PP5[7]);
  UBFA_8 U7 (W0[9], W2[8], PP0[8], PP1[8], PP2[8]);
  UBFA_8 U8 (W1[9], W3[8], PP3[8], PP4[8], PP5[8]);
  UBFA_9 U9 (W0[10], W2[9], PP0[9], PP1[9], PP2[9]);
  UBFA_9 U10 (W1[10], W3[9], PP3[9], PP4[9], PP5[9]);
  UBFA_10 U11 (W0[11], W2[10], PP0[10], PP1[10], PP2[10]);
  UBFA_10 U12 (W1[11], W3[10], PP3[10], PP4[10], PP5[10]);
  UBFA_11 U13 (W0[12], W2[11], PP0[11], PP1[11], PP2[11]);
  UBFA_11 U14 (W1[12], W3[11], PP3[11], PP4[11], PP5[11]);
  UBFA_12 U15 (W0[13], W2[12], PP0[12], PP1[12], PP2[12]);
  UBFA_12 U16 (W1[13], W3[12], PP3[12], PP4[12], PP5[12]);
  UBFA_13 U17 (W0[14], W2[13], PP0[13], PP1[13], PP2[13]);
  UBFA_13 U18 (W1[14], W3[13], PP3[13], PP4[13], PP5[13]);
  UBFA_14 U19 (W0[15], W2[14], PP0[14], PP1[14], PP2[14]);
  UBFA_14 U20 (W1[15], W3[14], PP3[14], PP4[14], PP5[14]);
  UBFA_15 U21 (W0[16], W2[15], PP0[15], PP1[15], PP2[15]);
  UBFA_15 U22 (W1[16], W3[15], PP3[15], PP4[15], PP5[15]);
  UBFA_16 U23 (W0[17], W2[16], PP0[16], PP1[16], PP2[16]);
  UBFA_16 U24 (W1[17], W3[16], PP3[16], PP4[16], PP5[16]);
  UBFA_17 U25 (W0[18], W2[17], PP0[17], PP1[17], PP2[17]);
  UBFA_17 U26 (W1[18], W3[17], PP3[17], PP4[17], PP5[17]);
  UBFA_18 U27 (W0[19], W2[18], PP0[18], PP1[18], PP2[18]);
  UBFA_18 U28 (W1[19], W3[18], PP3[18], PP4[18], PP5[18]);
  UBFA_19 U29 (W0[20], W2[19], PP0[19], PP1[19], PP2[19]);
  UBFA_19 U30 (W1[20], W3[19], PP3[19], PP4[19], PP5[19]);
  UBFA_20 U31 (W0[21], W2[20], PP0[20], PP1[20], PP2[20]);
  UBFA_20 U32 (W1[21], W3[20], PP3[20], PP4[20], PP5[20]);
  UBFA_21 U33 (W0[22], W2[21], PP0[21], PP1[21], PP2[21]);
  UBFA_21 U34 (W1[22], W3[21], PP3[21], PP4[21], PP5[21]);
  UBFA_22 U35 (W1[23], W2[22], PP0[22], PP1[22], PP2[22]);
  UBFA_22 U36 (W2[23], W3[22], PP3[22], PP4[22], PP5[22]);
  UBFA_23 U37 (W3[24], W3[23], PP0[23], PP1[23], PP2[23]);
  UBCON_3_0 U38 (W0[3:0], PP0[3:0]);
  UB1DCON_4 U39 (W0[4], PP2[4]);
  UB1DCON_5 U40 (W0[5], PP5[5]);
  UB1DCON_23 U41 (W0[23], PP3[23]);
  UBCON_26_24 U42 (W0[26:24], PP0[26:24]);
  UBCON_3_1 U43 (W1[3:1], PP1[3:1]);
  UB1DCON_4 U44 (W1[4], PP3[4]);
  UBCON_25_24 U45 (W1[25:24], PP1[25:24]);
  UBCON_3_2 U46 (W2[3:2], PP2[3:2]);
  UB1DCON_4 U47 (W2[4], PP4[4]);
  UB1DCON_24 U48 (W2[24], PP2[24]);
  UB1DCON_3 U49 (W3[3], PP3[3]);
  DADTR_26_0_25_1_2003 U50 (S1, S2, W0, W1, W2, W3);
endmodule

module DADTR_26_0_25_1_2003 (S1, S2, PP0, PP1, PP2, PP3);
  output [26:0] S1;
  output [26:1] S2;
  input [26:0] PP0;
  input [25:1] PP1;
  input [24:2] PP2;
  input [24:3] PP3;
  wire [26:0] W0;
  wire [25:1] W1;
  wire [25:2] W2;
  UBHA_3 U0 (W1[4], W2[3], PP0[3], PP1[3]);
  UBFA_4 U1 (W1[5], W2[4], PP0[4], PP1[4], PP2[4]);
  UBFA_5 U2 (W1[6], W2[5], PP0[5], PP1[5], PP2[5]);
  UBFA_6 U3 (W1[7], W2[6], PP0[6], PP1[6], PP2[6]);
  UBFA_7 U4 (W1[8], W2[7], PP0[7], PP1[7], PP2[7]);
  UBFA_8 U5 (W1[9], W2[8], PP0[8], PP1[8], PP2[8]);
  UBFA_9 U6 (W1[10], W2[9], PP0[9], PP1[9], PP2[9]);
  UBFA_10 U7 (W1[11], W2[10], PP0[10], PP1[10], PP2[10]);
  UBFA_11 U8 (W1[12], W2[11], PP0[11], PP1[11], PP2[11]);
  UBFA_12 U9 (W1[13], W2[12], PP0[12], PP1[12], PP2[12]);
  UBFA_13 U10 (W1[14], W2[13], PP0[13], PP1[13], PP2[13]);
  UBFA_14 U11 (W1[15], W2[14], PP0[14], PP1[14], PP2[14]);
  UBFA_15 U12 (W1[16], W2[15], PP0[15], PP1[15], PP2[15]);
  UBFA_16 U13 (W1[17], W2[16], PP0[16], PP1[16], PP2[16]);
  UBFA_17 U14 (W1[18], W2[17], PP0[17], PP1[17], PP2[17]);
  UBFA_18 U15 (W1[19], W2[18], PP0[18], PP1[18], PP2[18]);
  UBFA_19 U16 (W1[20], W2[19], PP0[19], PP1[19], PP2[19]);
  UBFA_20 U17 (W1[21], W2[20], PP0[20], PP1[20], PP2[20]);
  UBFA_21 U18 (W1[22], W2[21], PP0[21], PP1[21], PP2[21]);
  UBFA_22 U19 (W1[23], W2[22], PP0[22], PP1[22], PP2[22]);
  UBFA_23 U20 (W1[24], W2[23], PP0[23], PP1[23], PP2[23]);
  UBFA_24 U21 (W2[25], W2[24], PP0[24], PP1[24], PP2[24]);
  UBCON_2_0 U22 (W0[2:0], PP0[2:0]);
  UB1DCON_3 U23 (W0[3], PP2[3]);
  UBCON_24_4 U24 (W0[24:4], PP3[24:4]);
  UBCON_26_25 U25 (W0[26:25], PP0[26:25]);
  UBCON_2_1 U26 (W1[2:1], PP1[2:1]);
  UB1DCON_3 U27 (W1[3], PP3[3]);
  UB1DCON_25 U28 (W1[25], PP1[25]);
  UB1DCON_2 U29 (W2[2], PP2[2]);
  DADTR_26_0_25_1_2004 U30 (S1, S2, W0, W1, W2);
endmodule

module DADTR_26_0_25_1_2004 (S1, S2, PP0, PP1, PP2);
  output [26:0] S1;
  output [26:1] S2;
  input [26:0] PP0;
  input [25:1] PP1;
  input [25:2] PP2;
  wire [26:0] W0;
  wire [26:1] W1;
  UBHA_2 U0 (W0[3], W1[2], PP0[2], PP1[2]);
  UBFA_3 U1 (W0[4], W1[3], PP0[3], PP1[3], PP2[3]);
  UBFA_4 U2 (W0[5], W1[4], PP0[4], PP1[4], PP2[4]);
  UBFA_5 U3 (W0[6], W1[5], PP0[5], PP1[5], PP2[5]);
  UBFA_6 U4 (W0[7], W1[6], PP0[6], PP1[6], PP2[6]);
  UBFA_7 U5 (W0[8], W1[7], PP0[7], PP1[7], PP2[7]);
  UBFA_8 U6 (W0[9], W1[8], PP0[8], PP1[8], PP2[8]);
  UBFA_9 U7 (W0[10], W1[9], PP0[9], PP1[9], PP2[9]);
  UBFA_10 U8 (W0[11], W1[10], PP0[10], PP1[10], PP2[10]);
  UBFA_11 U9 (W0[12], W1[11], PP0[11], PP1[11], PP2[11]);
  UBFA_12 U10 (W0[13], W1[12], PP0[12], PP1[12], PP2[12]);
  UBFA_13 U11 (W0[14], W1[13], PP0[13], PP1[13], PP2[13]);
  UBFA_14 U12 (W0[15], W1[14], PP0[14], PP1[14], PP2[14]);
  UBFA_15 U13 (W0[16], W1[15], PP0[15], PP1[15], PP2[15]);
  UBFA_16 U14 (W0[17], W1[16], PP0[16], PP1[16], PP2[16]);
  UBFA_17 U15 (W0[18], W1[17], PP0[17], PP1[17], PP2[17]);
  UBFA_18 U16 (W0[19], W1[18], PP0[18], PP1[18], PP2[18]);
  UBFA_19 U17 (W0[20], W1[19], PP0[19], PP1[19], PP2[19]);
  UBFA_20 U18 (W0[21], W1[20], PP0[20], PP1[20], PP2[20]);
  UBFA_21 U19 (W0[22], W1[21], PP0[21], PP1[21], PP2[21]);
  UBFA_22 U20 (W0[23], W1[22], PP0[22], PP1[22], PP2[22]);
  UBFA_23 U21 (W0[24], W1[23], PP0[23], PP1[23], PP2[23]);
  UBFA_24 U22 (W0[25], W1[24], PP0[24], PP1[24], PP2[24]);
  UBFA_25 U23 (W1[26], W1[25], PP0[25], PP1[25], PP2[25]);
  UBCON_1_0 U24 (W0[1:0], PP0[1:0]);
  UB1DCON_2 U25 (W0[2], PP2[2]);
  UB1DCON_26 U26 (W0[26], PP0[26]);
  UB1DCON_1 U27 (W1[1], PP1[1]);
  DADTR_26_0_26_1 U28 (S1, S2, W0, W1);
endmodule

module DADTR_26_0_26_1 (S1, S2, PP0, PP1);
  output [26:0] S1;
  output [26:1] S2;
  input [26:0] PP0;
  input [26:1] PP1;
  UBCON_26_0 U0 (S1, PP0);
  UBCON_26_1 U1 (S2, PP1);
endmodule

module MultUB_STD_DAD_BC000 (P, IN1, IN2);
  output [27:0] P;
  input [13:0] IN1;
  input [13:0] IN2;
  wire [13:0] PP0;
  wire [14:1] PP1;
  wire [23:10] PP10;
  wire [24:11] PP11;
  wire [25:12] PP12;
  wire [26:13] PP13;
  wire [15:2] PP2;
  wire [16:3] PP3;
  wire [17:4] PP4;
  wire [18:5] PP5;
  wire [19:6] PP6;
  wire [20:7] PP7;
  wire [21:8] PP8;
  wire [22:9] PP9;
  wire [26:0] S1;
  wire [26:1] S2;
  UBPPG_13_0_13_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, IN1, IN2);
  DADTR_13_0_14_1_1000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13);
  UBBCL_26_0_26_1 U2 (P, S1, S2);
endmodule

module UBBCL_26_0_26_1 (S, X, Y);
  output [27:0] S;
  input [26:0] X;
  input [26:1] Y;
  UBPureBCL_26_1 U0 (S[27:1], X[26:1], Y[26:1]);
  UB1DCON_0 U1 (S[0], X[0]);
endmodule

module UBCON_12_0 (O, I);
  output [12:0] O;
  input [12:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
endmodule

module UBCON_12_1 (O, I);
  output [12:1] O;
  input [12:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
  UB1DCON_6 U5 (O[6], I[6]);
  UB1DCON_7 U6 (O[7], I[7]);
  UB1DCON_8 U7 (O[8], I[8]);
  UB1DCON_9 U8 (O[9], I[9]);
  UB1DCON_10 U9 (O[10], I[10]);
  UB1DCON_11 U10 (O[11], I[11]);
  UB1DCON_12 U11 (O[12], I[12]);
endmodule

module UBCON_12_10 (O, I);
  output [12:10] O;
  input [12:10] I;
  UB1DCON_10 U0 (O[10], I[10]);
  UB1DCON_11 U1 (O[11], I[11]);
  UB1DCON_12 U2 (O[12], I[12]);
endmodule

module UBCON_12_11 (O, I);
  output [12:11] O;
  input [12:11] I;
  UB1DCON_11 U0 (O[11], I[11]);
  UB1DCON_12 U1 (O[12], I[12]);
endmodule

module UBCON_12_2 (O, I);
  output [12:2] O;
  input [12:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
  UB1DCON_6 U4 (O[6], I[6]);
  UB1DCON_7 U5 (O[7], I[7]);
  UB1DCON_8 U6 (O[8], I[8]);
  UB1DCON_9 U7 (O[9], I[9]);
  UB1DCON_10 U8 (O[10], I[10]);
  UB1DCON_11 U9 (O[11], I[11]);
  UB1DCON_12 U10 (O[12], I[12]);
endmodule

module UBCON_12_3 (O, I);
  output [12:3] O;
  input [12:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
  UB1DCON_6 U3 (O[6], I[6]);
  UB1DCON_7 U4 (O[7], I[7]);
  UB1DCON_8 U5 (O[8], I[8]);
  UB1DCON_9 U6 (O[9], I[9]);
  UB1DCON_10 U7 (O[10], I[10]);
  UB1DCON_11 U8 (O[11], I[11]);
  UB1DCON_12 U9 (O[12], I[12]);
endmodule

module UBCON_12_4 (O, I);
  output [12:4] O;
  input [12:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
  UB1DCON_11 U7 (O[11], I[11]);
  UB1DCON_12 U8 (O[12], I[12]);
endmodule

module UBCON_12_5 (O, I);
  output [12:5] O;
  input [12:5] I;
  UB1DCON_5 U0 (O[5], I[5]);
  UB1DCON_6 U1 (O[6], I[6]);
  UB1DCON_7 U2 (O[7], I[7]);
  UB1DCON_8 U3 (O[8], I[8]);
  UB1DCON_9 U4 (O[9], I[9]);
  UB1DCON_10 U5 (O[10], I[10]);
  UB1DCON_11 U6 (O[11], I[11]);
  UB1DCON_12 U7 (O[12], I[12]);
endmodule

module UBCON_12_6 (O, I);
  output [12:6] O;
  input [12:6] I;
  UB1DCON_6 U0 (O[6], I[6]);
  UB1DCON_7 U1 (O[7], I[7]);
  UB1DCON_8 U2 (O[8], I[8]);
  UB1DCON_9 U3 (O[9], I[9]);
  UB1DCON_10 U4 (O[10], I[10]);
  UB1DCON_11 U5 (O[11], I[11]);
  UB1DCON_12 U6 (O[12], I[12]);
endmodule

module UBCON_12_7 (O, I);
  output [12:7] O;
  input [12:7] I;
  UB1DCON_7 U0 (O[7], I[7]);
  UB1DCON_8 U1 (O[8], I[8]);
  UB1DCON_9 U2 (O[9], I[9]);
  UB1DCON_10 U3 (O[10], I[10]);
  UB1DCON_11 U4 (O[11], I[11]);
  UB1DCON_12 U5 (O[12], I[12]);
endmodule

module UBCON_12_8 (O, I);
  output [12:8] O;
  input [12:8] I;
  UB1DCON_8 U0 (O[8], I[8]);
  UB1DCON_9 U1 (O[9], I[9]);
  UB1DCON_10 U2 (O[10], I[10]);
  UB1DCON_11 U3 (O[11], I[11]);
  UB1DCON_12 U4 (O[12], I[12]);
endmodule

module UBCON_12_9 (O, I);
  output [12:9] O;
  input [12:9] I;
  UB1DCON_9 U0 (O[9], I[9]);
  UB1DCON_10 U1 (O[10], I[10]);
  UB1DCON_11 U2 (O[11], I[11]);
  UB1DCON_12 U3 (O[12], I[12]);
endmodule

module UBCON_15_13 (O, I);
  output [15:13] O;
  input [15:13] I;
  UB1DCON_13 U0 (O[13], I[13]);
  UB1DCON_14 U1 (O[14], I[14]);
  UB1DCON_15 U2 (O[15], I[15]);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_20_19 (O, I);
  output [20:19] O;
  input [20:19] I;
  UB1DCON_19 U0 (O[19], I[19]);
  UB1DCON_20 U1 (O[20], I[20]);
endmodule

module UBCON_21_19 (O, I);
  output [21:19] O;
  input [21:19] I;
  UB1DCON_19 U0 (O[19], I[19]);
  UB1DCON_20 U1 (O[20], I[20]);
  UB1DCON_21 U2 (O[21], I[21]);
endmodule

module UBCON_22_19 (O, I);
  output [22:19] O;
  input [22:19] I;
  UB1DCON_19 U0 (O[19], I[19]);
  UB1DCON_20 U1 (O[20], I[20]);
  UB1DCON_21 U2 (O[21], I[21]);
  UB1DCON_22 U3 (O[22], I[22]);
endmodule

module UBCON_23_19 (O, I);
  output [23:19] O;
  input [23:19] I;
  UB1DCON_19 U0 (O[19], I[19]);
  UB1DCON_20 U1 (O[20], I[20]);
  UB1DCON_21 U2 (O[21], I[21]);
  UB1DCON_22 U3 (O[22], I[22]);
  UB1DCON_23 U4 (O[23], I[23]);
endmodule

module UBCON_23_22 (O, I);
  output [23:22] O;
  input [23:22] I;
  UB1DCON_22 U0 (O[22], I[22]);
  UB1DCON_23 U1 (O[23], I[23]);
endmodule

module UBCON_24_19 (O, I);
  output [24:19] O;
  input [24:19] I;
  UB1DCON_19 U0 (O[19], I[19]);
  UB1DCON_20 U1 (O[20], I[20]);
  UB1DCON_21 U2 (O[21], I[21]);
  UB1DCON_22 U3 (O[22], I[22]);
  UB1DCON_23 U4 (O[23], I[23]);
  UB1DCON_24 U5 (O[24], I[24]);
endmodule

module UBCON_24_22 (O, I);
  output [24:22] O;
  input [24:22] I;
  UB1DCON_22 U0 (O[22], I[22]);
  UB1DCON_23 U1 (O[23], I[23]);
  UB1DCON_24 U2 (O[24], I[24]);
endmodule

module UBCON_24_4 (O, I);
  output [24:4] O;
  input [24:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
  UB1DCON_11 U7 (O[11], I[11]);
  UB1DCON_12 U8 (O[12], I[12]);
  UB1DCON_13 U9 (O[13], I[13]);
  UB1DCON_14 U10 (O[14], I[14]);
  UB1DCON_15 U11 (O[15], I[15]);
  UB1DCON_16 U12 (O[16], I[16]);
  UB1DCON_17 U13 (O[17], I[17]);
  UB1DCON_18 U14 (O[18], I[18]);
  UB1DCON_19 U15 (O[19], I[19]);
  UB1DCON_20 U16 (O[20], I[20]);
  UB1DCON_21 U17 (O[21], I[21]);
  UB1DCON_22 U18 (O[22], I[22]);
  UB1DCON_23 U19 (O[23], I[23]);
  UB1DCON_24 U20 (O[24], I[24]);
endmodule

module UBCON_25_19 (O, I);
  output [25:19] O;
  input [25:19] I;
  UB1DCON_19 U0 (O[19], I[19]);
  UB1DCON_20 U1 (O[20], I[20]);
  UB1DCON_21 U2 (O[21], I[21]);
  UB1DCON_22 U3 (O[22], I[22]);
  UB1DCON_23 U4 (O[23], I[23]);
  UB1DCON_24 U5 (O[24], I[24]);
  UB1DCON_25 U6 (O[25], I[25]);
endmodule

module UBCON_25_22 (O, I);
  output [25:22] O;
  input [25:22] I;
  UB1DCON_22 U0 (O[22], I[22]);
  UB1DCON_23 U1 (O[23], I[23]);
  UB1DCON_24 U2 (O[24], I[24]);
  UB1DCON_25 U3 (O[25], I[25]);
endmodule

module UBCON_25_24 (O, I);
  output [25:24] O;
  input [25:24] I;
  UB1DCON_24 U0 (O[24], I[24]);
  UB1DCON_25 U1 (O[25], I[25]);
endmodule

module UBCON_26_0 (O, I);
  output [26:0] O;
  input [26:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
  UB1DCON_13 U13 (O[13], I[13]);
  UB1DCON_14 U14 (O[14], I[14]);
  UB1DCON_15 U15 (O[15], I[15]);
  UB1DCON_16 U16 (O[16], I[16]);
  UB1DCON_17 U17 (O[17], I[17]);
  UB1DCON_18 U18 (O[18], I[18]);
  UB1DCON_19 U19 (O[19], I[19]);
  UB1DCON_20 U20 (O[20], I[20]);
  UB1DCON_21 U21 (O[21], I[21]);
  UB1DCON_22 U22 (O[22], I[22]);
  UB1DCON_23 U23 (O[23], I[23]);
  UB1DCON_24 U24 (O[24], I[24]);
  UB1DCON_25 U25 (O[25], I[25]);
  UB1DCON_26 U26 (O[26], I[26]);
endmodule

module UBCON_26_1 (O, I);
  output [26:1] O;
  input [26:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
  UB1DCON_6 U5 (O[6], I[6]);
  UB1DCON_7 U6 (O[7], I[7]);
  UB1DCON_8 U7 (O[8], I[8]);
  UB1DCON_9 U8 (O[9], I[9]);
  UB1DCON_10 U9 (O[10], I[10]);
  UB1DCON_11 U10 (O[11], I[11]);
  UB1DCON_12 U11 (O[12], I[12]);
  UB1DCON_13 U12 (O[13], I[13]);
  UB1DCON_14 U13 (O[14], I[14]);
  UB1DCON_15 U14 (O[15], I[15]);
  UB1DCON_16 U15 (O[16], I[16]);
  UB1DCON_17 U16 (O[17], I[17]);
  UB1DCON_18 U17 (O[18], I[18]);
  UB1DCON_19 U18 (O[19], I[19]);
  UB1DCON_20 U19 (O[20], I[20]);
  UB1DCON_21 U20 (O[21], I[21]);
  UB1DCON_22 U21 (O[22], I[22]);
  UB1DCON_23 U22 (O[23], I[23]);
  UB1DCON_24 U23 (O[24], I[24]);
  UB1DCON_25 U24 (O[25], I[25]);
  UB1DCON_26 U25 (O[26], I[26]);
endmodule

module UBCON_26_19 (O, I);
  output [26:19] O;
  input [26:19] I;
  UB1DCON_19 U0 (O[19], I[19]);
  UB1DCON_20 U1 (O[20], I[20]);
  UB1DCON_21 U2 (O[21], I[21]);
  UB1DCON_22 U3 (O[22], I[22]);
  UB1DCON_23 U4 (O[23], I[23]);
  UB1DCON_24 U5 (O[24], I[24]);
  UB1DCON_25 U6 (O[25], I[25]);
  UB1DCON_26 U7 (O[26], I[26]);
endmodule

module UBCON_26_22 (O, I);
  output [26:22] O;
  input [26:22] I;
  UB1DCON_22 U0 (O[22], I[22]);
  UB1DCON_23 U1 (O[23], I[23]);
  UB1DCON_24 U2 (O[24], I[24]);
  UB1DCON_25 U3 (O[25], I[25]);
  UB1DCON_26 U4 (O[26], I[26]);
endmodule

module UBCON_26_24 (O, I);
  output [26:24] O;
  input [26:24] I;
  UB1DCON_24 U0 (O[24], I[24]);
  UB1DCON_25 U1 (O[25], I[25]);
  UB1DCON_26 U2 (O[26], I[26]);
endmodule

module UBCON_26_25 (O, I);
  output [26:25] O;
  input [26:25] I;
  UB1DCON_25 U0 (O[25], I[25]);
  UB1DCON_26 U1 (O[26], I[26]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBCON_2_1 (O, I);
  output [2:1] O;
  input [2:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
endmodule

module UBCON_3_0 (O, I);
  output [3:0] O;
  input [3:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
endmodule

module UBCON_3_1 (O, I);
  output [3:1] O;
  input [3:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
endmodule

module UBCON_3_2 (O, I);
  output [3:2] O;
  input [3:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
endmodule

module UBCON_5_0 (O, I);
  output [5:0] O;
  input [5:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
endmodule

module UBCON_5_1 (O, I);
  output [5:1] O;
  input [5:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
endmodule

module UBCON_5_2 (O, I);
  output [5:2] O;
  input [5:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
endmodule

module UBCON_5_3 (O, I);
  output [5:3] O;
  input [5:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
endmodule

module UBCON_5_4 (O, I);
  output [5:4] O;
  input [5:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
endmodule

module UBCON_8_0 (O, I);
  output [8:0] O;
  input [8:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
endmodule

module UBCON_8_1 (O, I);
  output [8:1] O;
  input [8:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
  UB1DCON_6 U5 (O[6], I[6]);
  UB1DCON_7 U6 (O[7], I[7]);
  UB1DCON_8 U7 (O[8], I[8]);
endmodule

module UBCON_8_2 (O, I);
  output [8:2] O;
  input [8:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
  UB1DCON_6 U4 (O[6], I[6]);
  UB1DCON_7 U5 (O[7], I[7]);
  UB1DCON_8 U6 (O[8], I[8]);
endmodule

module UBCON_8_3 (O, I);
  output [8:3] O;
  input [8:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
  UB1DCON_6 U3 (O[6], I[6]);
  UB1DCON_7 U4 (O[7], I[7]);
  UB1DCON_8 U5 (O[8], I[8]);
endmodule

module UBCON_8_4 (O, I);
  output [8:4] O;
  input [8:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
endmodule

module UBCON_8_5 (O, I);
  output [8:5] O;
  input [8:5] I;
  UB1DCON_5 U0 (O[5], I[5]);
  UB1DCON_6 U1 (O[6], I[6]);
  UB1DCON_7 U2 (O[7], I[7]);
  UB1DCON_8 U3 (O[8], I[8]);
endmodule

module UBCON_8_6 (O, I);
  output [8:6] O;
  input [8:6] I;
  UB1DCON_6 U0 (O[6], I[6]);
  UB1DCON_7 U1 (O[7], I[7]);
  UB1DCON_8 U2 (O[8], I[8]);
endmodule

module UBCON_8_7 (O, I);
  output [8:7] O;
  input [8:7] I;
  UB1DCON_7 U0 (O[7], I[7]);
  UB1DCON_8 U1 (O[8], I[8]);
endmodule

module UBPPG_13_0_13_0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, IN1, IN2);
  output [13:0] PP0;
  output [14:1] PP1;
  output [23:10] PP10;
  output [24:11] PP11;
  output [25:12] PP12;
  output [26:13] PP13;
  output [15:2] PP2;
  output [16:3] PP3;
  output [17:4] PP4;
  output [18:5] PP5;
  output [19:6] PP6;
  output [20:7] PP7;
  output [21:8] PP8;
  output [22:9] PP9;
  input [13:0] IN1;
  input [13:0] IN2;
  UBVPPG_13_0_0 U0 (PP0, IN1, IN2[0]);
  UBVPPG_13_0_1 U1 (PP1, IN1, IN2[1]);
  UBVPPG_13_0_2 U2 (PP2, IN1, IN2[2]);
  UBVPPG_13_0_3 U3 (PP3, IN1, IN2[3]);
  UBVPPG_13_0_4 U4 (PP4, IN1, IN2[4]);
  UBVPPG_13_0_5 U5 (PP5, IN1, IN2[5]);
  UBVPPG_13_0_6 U6 (PP6, IN1, IN2[6]);
  UBVPPG_13_0_7 U7 (PP7, IN1, IN2[7]);
  UBVPPG_13_0_8 U8 (PP8, IN1, IN2[8]);
  UBVPPG_13_0_9 U9 (PP9, IN1, IN2[9]);
  UBVPPG_13_0_10 U10 (PP10, IN1, IN2[10]);
  UBVPPG_13_0_11 U11 (PP11, IN1, IN2[11]);
  UBVPPG_13_0_12 U12 (PP12, IN1, IN2[12]);
  UBVPPG_13_0_13 U13 (PP13, IN1, IN2[13]);
endmodule

module UBPureBCL_26_1 (S, X, Y);
  output [27:1] S;
  input [26:1] X;
  input [26:1] Y;
  wire C;
  PriMBCLA_26_1 U0 (S, X, Y, C);
  UBZero_1_1 U1 (C);
endmodule

module UBVPPG_13_0_0 (O, IN1, IN2);
  output [13:0] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
  UB1BPPG_6_0 U6 (O[6], IN1[6], IN2);
  UB1BPPG_7_0 U7 (O[7], IN1[7], IN2);
  UB1BPPG_8_0 U8 (O[8], IN1[8], IN2);
  UB1BPPG_9_0 U9 (O[9], IN1[9], IN2);
  UB1BPPG_10_0 U10 (O[10], IN1[10], IN2);
  UB1BPPG_11_0 U11 (O[11], IN1[11], IN2);
  UB1BPPG_12_0 U12 (O[12], IN1[12], IN2);
  UB1BPPG_13_0 U13 (O[13], IN1[13], IN2);
endmodule

module UBVPPG_13_0_1 (O, IN1, IN2);
  output [14:1] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_1 U0 (O[1], IN1[0], IN2);
  UB1BPPG_1_1 U1 (O[2], IN1[1], IN2);
  UB1BPPG_2_1 U2 (O[3], IN1[2], IN2);
  UB1BPPG_3_1 U3 (O[4], IN1[3], IN2);
  UB1BPPG_4_1 U4 (O[5], IN1[4], IN2);
  UB1BPPG_5_1 U5 (O[6], IN1[5], IN2);
  UB1BPPG_6_1 U6 (O[7], IN1[6], IN2);
  UB1BPPG_7_1 U7 (O[8], IN1[7], IN2);
  UB1BPPG_8_1 U8 (O[9], IN1[8], IN2);
  UB1BPPG_9_1 U9 (O[10], IN1[9], IN2);
  UB1BPPG_10_1 U10 (O[11], IN1[10], IN2);
  UB1BPPG_11_1 U11 (O[12], IN1[11], IN2);
  UB1BPPG_12_1 U12 (O[13], IN1[12], IN2);
  UB1BPPG_13_1 U13 (O[14], IN1[13], IN2);
endmodule

module UBVPPG_13_0_10 (O, IN1, IN2);
  output [23:10] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_10 U0 (O[10], IN1[0], IN2);
  UB1BPPG_1_10 U1 (O[11], IN1[1], IN2);
  UB1BPPG_2_10 U2 (O[12], IN1[2], IN2);
  UB1BPPG_3_10 U3 (O[13], IN1[3], IN2);
  UB1BPPG_4_10 U4 (O[14], IN1[4], IN2);
  UB1BPPG_5_10 U5 (O[15], IN1[5], IN2);
  UB1BPPG_6_10 U6 (O[16], IN1[6], IN2);
  UB1BPPG_7_10 U7 (O[17], IN1[7], IN2);
  UB1BPPG_8_10 U8 (O[18], IN1[8], IN2);
  UB1BPPG_9_10 U9 (O[19], IN1[9], IN2);
  UB1BPPG_10_10 U10 (O[20], IN1[10], IN2);
  UB1BPPG_11_10 U11 (O[21], IN1[11], IN2);
  UB1BPPG_12_10 U12 (O[22], IN1[12], IN2);
  UB1BPPG_13_10 U13 (O[23], IN1[13], IN2);
endmodule

module UBVPPG_13_0_11 (O, IN1, IN2);
  output [24:11] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_11 U0 (O[11], IN1[0], IN2);
  UB1BPPG_1_11 U1 (O[12], IN1[1], IN2);
  UB1BPPG_2_11 U2 (O[13], IN1[2], IN2);
  UB1BPPG_3_11 U3 (O[14], IN1[3], IN2);
  UB1BPPG_4_11 U4 (O[15], IN1[4], IN2);
  UB1BPPG_5_11 U5 (O[16], IN1[5], IN2);
  UB1BPPG_6_11 U6 (O[17], IN1[6], IN2);
  UB1BPPG_7_11 U7 (O[18], IN1[7], IN2);
  UB1BPPG_8_11 U8 (O[19], IN1[8], IN2);
  UB1BPPG_9_11 U9 (O[20], IN1[9], IN2);
  UB1BPPG_10_11 U10 (O[21], IN1[10], IN2);
  UB1BPPG_11_11 U11 (O[22], IN1[11], IN2);
  UB1BPPG_12_11 U12 (O[23], IN1[12], IN2);
  UB1BPPG_13_11 U13 (O[24], IN1[13], IN2);
endmodule

module UBVPPG_13_0_12 (O, IN1, IN2);
  output [25:12] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_12 U0 (O[12], IN1[0], IN2);
  UB1BPPG_1_12 U1 (O[13], IN1[1], IN2);
  UB1BPPG_2_12 U2 (O[14], IN1[2], IN2);
  UB1BPPG_3_12 U3 (O[15], IN1[3], IN2);
  UB1BPPG_4_12 U4 (O[16], IN1[4], IN2);
  UB1BPPG_5_12 U5 (O[17], IN1[5], IN2);
  UB1BPPG_6_12 U6 (O[18], IN1[6], IN2);
  UB1BPPG_7_12 U7 (O[19], IN1[7], IN2);
  UB1BPPG_8_12 U8 (O[20], IN1[8], IN2);
  UB1BPPG_9_12 U9 (O[21], IN1[9], IN2);
  UB1BPPG_10_12 U10 (O[22], IN1[10], IN2);
  UB1BPPG_11_12 U11 (O[23], IN1[11], IN2);
  UB1BPPG_12_12 U12 (O[24], IN1[12], IN2);
  UB1BPPG_13_12 U13 (O[25], IN1[13], IN2);
endmodule

module UBVPPG_13_0_13 (O, IN1, IN2);
  output [26:13] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_13 U0 (O[13], IN1[0], IN2);
  UB1BPPG_1_13 U1 (O[14], IN1[1], IN2);
  UB1BPPG_2_13 U2 (O[15], IN1[2], IN2);
  UB1BPPG_3_13 U3 (O[16], IN1[3], IN2);
  UB1BPPG_4_13 U4 (O[17], IN1[4], IN2);
  UB1BPPG_5_13 U5 (O[18], IN1[5], IN2);
  UB1BPPG_6_13 U6 (O[19], IN1[6], IN2);
  UB1BPPG_7_13 U7 (O[20], IN1[7], IN2);
  UB1BPPG_8_13 U8 (O[21], IN1[8], IN2);
  UB1BPPG_9_13 U9 (O[22], IN1[9], IN2);
  UB1BPPG_10_13 U10 (O[23], IN1[10], IN2);
  UB1BPPG_11_13 U11 (O[24], IN1[11], IN2);
  UB1BPPG_12_13 U12 (O[25], IN1[12], IN2);
  UB1BPPG_13_13 U13 (O[26], IN1[13], IN2);
endmodule

module UBVPPG_13_0_2 (O, IN1, IN2);
  output [15:2] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
  UB1BPPG_6_2 U6 (O[8], IN1[6], IN2);
  UB1BPPG_7_2 U7 (O[9], IN1[7], IN2);
  UB1BPPG_8_2 U8 (O[10], IN1[8], IN2);
  UB1BPPG_9_2 U9 (O[11], IN1[9], IN2);
  UB1BPPG_10_2 U10 (O[12], IN1[10], IN2);
  UB1BPPG_11_2 U11 (O[13], IN1[11], IN2);
  UB1BPPG_12_2 U12 (O[14], IN1[12], IN2);
  UB1BPPG_13_2 U13 (O[15], IN1[13], IN2);
endmodule

module UBVPPG_13_0_3 (O, IN1, IN2);
  output [16:3] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_3 U0 (O[3], IN1[0], IN2);
  UB1BPPG_1_3 U1 (O[4], IN1[1], IN2);
  UB1BPPG_2_3 U2 (O[5], IN1[2], IN2);
  UB1BPPG_3_3 U3 (O[6], IN1[3], IN2);
  UB1BPPG_4_3 U4 (O[7], IN1[4], IN2);
  UB1BPPG_5_3 U5 (O[8], IN1[5], IN2);
  UB1BPPG_6_3 U6 (O[9], IN1[6], IN2);
  UB1BPPG_7_3 U7 (O[10], IN1[7], IN2);
  UB1BPPG_8_3 U8 (O[11], IN1[8], IN2);
  UB1BPPG_9_3 U9 (O[12], IN1[9], IN2);
  UB1BPPG_10_3 U10 (O[13], IN1[10], IN2);
  UB1BPPG_11_3 U11 (O[14], IN1[11], IN2);
  UB1BPPG_12_3 U12 (O[15], IN1[12], IN2);
  UB1BPPG_13_3 U13 (O[16], IN1[13], IN2);
endmodule

module UBVPPG_13_0_4 (O, IN1, IN2);
  output [17:4] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
  UB1BPPG_6_4 U6 (O[10], IN1[6], IN2);
  UB1BPPG_7_4 U7 (O[11], IN1[7], IN2);
  UB1BPPG_8_4 U8 (O[12], IN1[8], IN2);
  UB1BPPG_9_4 U9 (O[13], IN1[9], IN2);
  UB1BPPG_10_4 U10 (O[14], IN1[10], IN2);
  UB1BPPG_11_4 U11 (O[15], IN1[11], IN2);
  UB1BPPG_12_4 U12 (O[16], IN1[12], IN2);
  UB1BPPG_13_4 U13 (O[17], IN1[13], IN2);
endmodule

module UBVPPG_13_0_5 (O, IN1, IN2);
  output [18:5] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_5 U0 (O[5], IN1[0], IN2);
  UB1BPPG_1_5 U1 (O[6], IN1[1], IN2);
  UB1BPPG_2_5 U2 (O[7], IN1[2], IN2);
  UB1BPPG_3_5 U3 (O[8], IN1[3], IN2);
  UB1BPPG_4_5 U4 (O[9], IN1[4], IN2);
  UB1BPPG_5_5 U5 (O[10], IN1[5], IN2);
  UB1BPPG_6_5 U6 (O[11], IN1[6], IN2);
  UB1BPPG_7_5 U7 (O[12], IN1[7], IN2);
  UB1BPPG_8_5 U8 (O[13], IN1[8], IN2);
  UB1BPPG_9_5 U9 (O[14], IN1[9], IN2);
  UB1BPPG_10_5 U10 (O[15], IN1[10], IN2);
  UB1BPPG_11_5 U11 (O[16], IN1[11], IN2);
  UB1BPPG_12_5 U12 (O[17], IN1[12], IN2);
  UB1BPPG_13_5 U13 (O[18], IN1[13], IN2);
endmodule

module UBVPPG_13_0_6 (O, IN1, IN2);
  output [19:6] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_6 U0 (O[6], IN1[0], IN2);
  UB1BPPG_1_6 U1 (O[7], IN1[1], IN2);
  UB1BPPG_2_6 U2 (O[8], IN1[2], IN2);
  UB1BPPG_3_6 U3 (O[9], IN1[3], IN2);
  UB1BPPG_4_6 U4 (O[10], IN1[4], IN2);
  UB1BPPG_5_6 U5 (O[11], IN1[5], IN2);
  UB1BPPG_6_6 U6 (O[12], IN1[6], IN2);
  UB1BPPG_7_6 U7 (O[13], IN1[7], IN2);
  UB1BPPG_8_6 U8 (O[14], IN1[8], IN2);
  UB1BPPG_9_6 U9 (O[15], IN1[9], IN2);
  UB1BPPG_10_6 U10 (O[16], IN1[10], IN2);
  UB1BPPG_11_6 U11 (O[17], IN1[11], IN2);
  UB1BPPG_12_6 U12 (O[18], IN1[12], IN2);
  UB1BPPG_13_6 U13 (O[19], IN1[13], IN2);
endmodule

module UBVPPG_13_0_7 (O, IN1, IN2);
  output [20:7] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_7 U0 (O[7], IN1[0], IN2);
  UB1BPPG_1_7 U1 (O[8], IN1[1], IN2);
  UB1BPPG_2_7 U2 (O[9], IN1[2], IN2);
  UB1BPPG_3_7 U3 (O[10], IN1[3], IN2);
  UB1BPPG_4_7 U4 (O[11], IN1[4], IN2);
  UB1BPPG_5_7 U5 (O[12], IN1[5], IN2);
  UB1BPPG_6_7 U6 (O[13], IN1[6], IN2);
  UB1BPPG_7_7 U7 (O[14], IN1[7], IN2);
  UB1BPPG_8_7 U8 (O[15], IN1[8], IN2);
  UB1BPPG_9_7 U9 (O[16], IN1[9], IN2);
  UB1BPPG_10_7 U10 (O[17], IN1[10], IN2);
  UB1BPPG_11_7 U11 (O[18], IN1[11], IN2);
  UB1BPPG_12_7 U12 (O[19], IN1[12], IN2);
  UB1BPPG_13_7 U13 (O[20], IN1[13], IN2);
endmodule

module UBVPPG_13_0_8 (O, IN1, IN2);
  output [21:8] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_8 U0 (O[8], IN1[0], IN2);
  UB1BPPG_1_8 U1 (O[9], IN1[1], IN2);
  UB1BPPG_2_8 U2 (O[10], IN1[2], IN2);
  UB1BPPG_3_8 U3 (O[11], IN1[3], IN2);
  UB1BPPG_4_8 U4 (O[12], IN1[4], IN2);
  UB1BPPG_5_8 U5 (O[13], IN1[5], IN2);
  UB1BPPG_6_8 U6 (O[14], IN1[6], IN2);
  UB1BPPG_7_8 U7 (O[15], IN1[7], IN2);
  UB1BPPG_8_8 U8 (O[16], IN1[8], IN2);
  UB1BPPG_9_8 U9 (O[17], IN1[9], IN2);
  UB1BPPG_10_8 U10 (O[18], IN1[10], IN2);
  UB1BPPG_11_8 U11 (O[19], IN1[11], IN2);
  UB1BPPG_12_8 U12 (O[20], IN1[12], IN2);
  UB1BPPG_13_8 U13 (O[21], IN1[13], IN2);
endmodule

module UBVPPG_13_0_9 (O, IN1, IN2);
  output [22:9] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_9 U0 (O[9], IN1[0], IN2);
  UB1BPPG_1_9 U1 (O[10], IN1[1], IN2);
  UB1BPPG_2_9 U2 (O[11], IN1[2], IN2);
  UB1BPPG_3_9 U3 (O[12], IN1[3], IN2);
  UB1BPPG_4_9 U4 (O[13], IN1[4], IN2);
  UB1BPPG_5_9 U5 (O[14], IN1[5], IN2);
  UB1BPPG_6_9 U6 (O[15], IN1[6], IN2);
  UB1BPPG_7_9 U7 (O[16], IN1[7], IN2);
  UB1BPPG_8_9 U8 (O[17], IN1[8], IN2);
  UB1BPPG_9_9 U9 (O[18], IN1[9], IN2);
  UB1BPPG_10_9 U10 (O[19], IN1[10], IN2);
  UB1BPPG_11_9 U11 (O[20], IN1[11], IN2);
  UB1BPPG_12_9 U12 (O[21], IN1[12], IN2);
  UB1BPPG_13_9 U13 (O[22], IN1[13], IN2);
endmodule

