/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: Multiplier_15_0_1000

  Number system: Unsigned binary
  Multiplicand length: 16
  Multiplier length: 16
  Partial product generation: Simple PPG
  Partial product accumulation: (4;2) compressor tree
  Final stage addition: Conditional sum adder
----------------------------------------------------------------------------*/

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_1(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_2(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBZero_3_3(O);
  output [3:3] O;
  assign O[3] = 0;
endmodule

module UB1B4_2CMP_3(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_4(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_5(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_6(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_7(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_8(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_9(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_10(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_11(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_12(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_13(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_14(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_15(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B3_2CMP_16(Co, C, S, IN0, IN1, IN2, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UBFA_17(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB1DCON_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_5(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBZero_7_7(O);
  output [7:7] O;
  assign O[7] = 0;
endmodule

module UB1B4_2CMP_16(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_17(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_18(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_19(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B3_2CMP_20(Co, C, S, IN0, IN1, IN2, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UBFA_21(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB1DCON_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_9(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBZero_11_11(O);
  output [11:11] O;
  assign O[11] = 0;
endmodule

module UB1B4_2CMP_20(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_21(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_22(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_23(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B3_2CMP_24(Co, C, S, IN0, IN1, IN2, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UBFA_25(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB1DCON_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_13(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_14(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBZero_15_15(O);
  output [15:15] O;
  assign O[15] = 0;
endmodule

module UB1B4_2CMP_24(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_25(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_26(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B4_2CMP_27(Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2 ^ IN3;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci ) | ( ~ W2 & IN3 );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UB1B3_2CMP_28(Co, C, S, IN0, IN1, IN2, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UBFA_29(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB1DCON_30(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBZero_6_6(O);
  output [6:6] O;
  assign O[6] = 0;
endmodule

module UBFA_19(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_20(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_21(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_22(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_10(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_11(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_12(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_13(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBZero_14_14(O);
  output [14:14] O;
  assign O[14] = 0;
endmodule

module UBFA_27(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_28(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_29(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_30(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_6(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_7(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB1B3_2CMP_23(Co, C, S, IN0, IN1, IN2, Ci);
  output C;
  output Co;
  output S;
  input Ci;
  input IN0;
  input IN1;
  input IN2;
  wire W0;
  wire W1;
  wire W2;
  assign W0 = IN0 ^ IN1;
  assign W1 = IN2;
  assign W2 = W0 ^ W1;
  assign S = W2 ^ Ci;
  assign C = ( W2 & Ci );
  assign Co = ( W0 & IN2 ) | ( ~ W0 & IN0 );
endmodule

module UBFA_24(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_25(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_26(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_27(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_31(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHCSuB_4_4(C, S, X, Y, Ci);
  output C;
  output S;
  input Ci;
  input X;
  input Y;
  UBFA_4 U0 (C, S, X, Y, Ci);
endmodule

module UBZero_5_5(O);
  output [5:5] O;
  assign O[5] = 0;
endmodule

module UBOne_5(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_5_5(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_5_5 U0 (Ci_0);
  UBOne_5 U1 (Ci_1);
  UBFA_5 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_5 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBHCSuB_5_4(C, S, X, Y, Ci);
  output C;
  output [5:4] S;
  input Ci;
  input [5:4] X;
  input [5:4] Y;
  wire C_0;
  wire C_1;
  wire Co;
  wire S_0;
  wire S_1;
  assign S[5] = ( S_0 & ( ~ Co ) ) | ( S_1 & Co );
  assign C = ( C_0 & ( ~ Co ) ) | ( C_1 & Co );
  UBHCSuB_4_4 U0 (Co, S[4], X[4], Y[4], Ci);
  UBCSuB_5_5 U1 (C_0, C_1, S_0, S_1, X[5], Y[5]);
endmodule

module UBOne_6(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_6_6(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_6_6 U0 (Ci_0);
  UBOne_6 U1 (Ci_1);
  UBFA_6 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_6 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_7(O);
  output O;
  assign O = 1;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSuB_7_7(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_7_7 U0 (Ci_0);
  UBOne_7 U1 (Ci_1);
  UBFA_7 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_7 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_7_6(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [7:6] S_0;
  output [7:6] S_1;
  input [7:6] X;
  input [7:6] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire So_0;
  wire So_1;
  assign S_0[7] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[7] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_6_6 U0 (Ci_0, Ci_1, S_0[6], S_1[6], X[6], Y[6]);
  UBCSuB_7_7 U1 (Co_0, Co_1, So_0, So_1, X[7], Y[7]);
endmodule

module UBHCSuB_7_4(C, S, X, Y, Ci);
  output C;
  output [7:4] S;
  input Ci;
  input [7:4] X;
  input [7:4] Y;
  wire C_0;
  wire C_1;
  wire Co;
  wire [7:6] S_0;
  wire [7:6] S_1;
  assign S[6] = ( S_0[6] & ( ~ Co ) ) | ( S_1[6] & Co );
  assign S[7] = ( S_0[7] & ( ~ Co ) ) | ( S_1[7] & Co );
  assign C = ( C_0 & ( ~ Co ) ) | ( C_1 & Co );
  UBHCSuB_5_4 U0 (Co, S[5:4], X[5:4], Y[5:4], Ci);
  UBCSuB_7_6 U1 (C_0, C_1, S_0, S_1, X[7:6], Y[7:6]);
endmodule

module UBZero_8_8(O);
  output [8:8] O;
  assign O[8] = 0;
endmodule

module UBOne_8(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_8_8(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_8_8 U0 (Ci_0);
  UBOne_8 U1 (Ci_1);
  UBFA_8 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_8 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBZero_9_9(O);
  output [9:9] O;
  assign O[9] = 0;
endmodule

module UBOne_9(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_9_9(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_9_9 U0 (Ci_0);
  UBOne_9 U1 (Ci_1);
  UBFA_9 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_9 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_9_8(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [9:8] S_0;
  output [9:8] S_1;
  input [9:8] X;
  input [9:8] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire So_0;
  wire So_1;
  assign S_0[9] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[9] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_8_8 U0 (Ci_0, Ci_1, S_0[8], S_1[8], X[8], Y[8]);
  UBCSuB_9_9 U1 (Co_0, Co_1, So_0, So_1, X[9], Y[9]);
endmodule

module UBZero_10_10(O);
  output [10:10] O;
  assign O[10] = 0;
endmodule

module UBOne_10(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_10_10(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_10_10 U0 (Ci_0);
  UBOne_10 U1 (Ci_1);
  UBFA_10 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_10 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_10_8(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [10:8] S_0;
  output [10:8] S_1;
  input [10:8] X;
  input [10:8] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [10:10] So_0;
  wire [10:10] So_1;
  assign S_0[10] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[10] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_9_8 U0 (Ci_0, Ci_1, S_0[9:8], S_1[9:8], X[9:8], Y[9:8]);
  UBCSuB_10_10 U1 (Co_0, Co_1, So_0, So_1, X[10], Y[10]);
endmodule

module UBHCSuB_10_4(C, S, X, Y, Ci);
  output C;
  output [10:4] S;
  input Ci;
  input [10:4] X;
  input [10:4] Y;
  wire C_0;
  wire C_1;
  wire Co;
  wire [10:8] S_0;
  wire [10:8] S_1;
  assign S[8] = ( S_0[8] & ( ~ Co ) ) | ( S_1[8] & Co );
  assign S[9] = ( S_0[9] & ( ~ Co ) ) | ( S_1[9] & Co );
  assign S[10] = ( S_0[10] & ( ~ Co ) ) | ( S_1[10] & Co );
  assign C = ( C_0 & ( ~ Co ) ) | ( C_1 & Co );
  UBHCSuB_7_4 U0 (Co, S[7:4], X[7:4], Y[7:4], Ci);
  UBCSuB_10_8 U1 (C_0, C_1, S_0, S_1, X[10:8], Y[10:8]);
endmodule

module UBOne_11(O);
  output O;
  assign O = 1;
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSuB_11_11(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_11_11 U0 (Ci_0);
  UBOne_11 U1 (Ci_1);
  UBFA_11 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_11 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBZero_12_12(O);
  output [12:12] O;
  assign O[12] = 0;
endmodule

module UBOne_12(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_12_12(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_12_12 U0 (Ci_0);
  UBOne_12 U1 (Ci_1);
  UBFA_12 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_12 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_12_11(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [12:11] S_0;
  output [12:11] S_1;
  input [12:11] X;
  input [12:11] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire So_0;
  wire So_1;
  assign S_0[12] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[12] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_11_11 U0 (Ci_0, Ci_1, S_0[11], S_1[11], X[11], Y[11]);
  UBCSuB_12_12 U1 (Co_0, Co_1, So_0, So_1, X[12], Y[12]);
endmodule

module UBZero_13_13(O);
  output [13:13] O;
  assign O[13] = 0;
endmodule

module UBOne_13(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_13_13(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_13_13 U0 (Ci_0);
  UBOne_13 U1 (Ci_1);
  UBFA_13 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_13 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_14(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_14_14(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_14_14 U0 (Ci_0);
  UBOne_14 U1 (Ci_1);
  UBFA_14 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_14 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_14_13(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [14:13] S_0;
  output [14:13] S_1;
  input [14:13] X;
  input [14:13] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire So_0;
  wire So_1;
  assign S_0[14] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[14] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_13_13 U0 (Ci_0, Ci_1, S_0[13], S_1[13], X[13], Y[13]);
  UBCSuB_14_14 U1 (Co_0, Co_1, So_0, So_1, X[14], Y[14]);
endmodule

module UBCSuB_14_11(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [14:11] S_0;
  output [14:11] S_1;
  input [14:11] X;
  input [14:11] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [14:13] So_0;
  wire [14:13] So_1;
  assign S_0[13] = ( So_0[13] & ( ~ Ci_0 ) ) | ( So_1[13] & Ci_0 );
  assign S_0[14] = ( So_0[14] & ( ~ Ci_0 ) ) | ( So_1[14] & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[13] = ( So_0[13] & ( ~ Ci_1 ) ) | ( So_1[13] & Ci_1 );
  assign S_1[14] = ( So_0[14] & ( ~ Ci_1 ) ) | ( So_1[14] & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_12_11 U0 (Ci_0, Ci_1, S_0[12:11], S_1[12:11], X[12:11], Y[12:11]);
  UBCSuB_14_13 U1 (Co_0, Co_1, So_0, So_1, X[14:13], Y[14:13]);
endmodule

module UBOne_15(O);
  output O;
  assign O = 1;
endmodule

module UBFA_15(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSuB_15_15(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_15_15 U0 (Ci_0);
  UBOne_15 U1 (Ci_1);
  UBFA_15 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_15 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBZero_16_16(O);
  output [16:16] O;
  assign O[16] = 0;
endmodule

module UBOne_16(O);
  output O;
  assign O = 1;
endmodule

module UBFA_16(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSuB_16_16(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_16_16 U0 (Ci_0);
  UBOne_16 U1 (Ci_1);
  UBFA_16 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_16 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_16_15(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [16:15] S_0;
  output [16:15] S_1;
  input [16:15] X;
  input [16:15] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire So_0;
  wire So_1;
  assign S_0[16] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[16] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_15_15 U0 (Ci_0, Ci_1, S_0[15], S_1[15], X[15], Y[15]);
  UBCSuB_16_16 U1 (Co_0, Co_1, So_0, So_1, X[16], Y[16]);
endmodule

module UBZero_17_17(O);
  output [17:17] O;
  assign O[17] = 0;
endmodule

module UBOne_17(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_17_17(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_17_17 U0 (Ci_0);
  UBOne_17 U1 (Ci_1);
  UBFA_17 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_17 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_17_15(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [17:15] S_0;
  output [17:15] S_1;
  input [17:15] X;
  input [17:15] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [17:17] So_0;
  wire [17:17] So_1;
  assign S_0[17] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[17] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_16_15 U0 (Ci_0, Ci_1, S_0[16:15], S_1[16:15], X[16:15], Y[16:15]);
  UBCSuB_17_17 U1 (Co_0, Co_1, So_0, So_1, X[17], Y[17]);
endmodule

module UBCSuB_17_11(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [17:11] S_0;
  output [17:11] S_1;
  input [17:11] X;
  input [17:11] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [17:15] So_0;
  wire [17:15] So_1;
  assign S_0[15] = ( So_0[15] & ( ~ Ci_0 ) ) | ( So_1[15] & Ci_0 );
  assign S_0[16] = ( So_0[16] & ( ~ Ci_0 ) ) | ( So_1[16] & Ci_0 );
  assign S_0[17] = ( So_0[17] & ( ~ Ci_0 ) ) | ( So_1[17] & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[15] = ( So_0[15] & ( ~ Ci_1 ) ) | ( So_1[15] & Ci_1 );
  assign S_1[16] = ( So_0[16] & ( ~ Ci_1 ) ) | ( So_1[16] & Ci_1 );
  assign S_1[17] = ( So_0[17] & ( ~ Ci_1 ) ) | ( So_1[17] & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_14_11 U0 (Ci_0, Ci_1, S_0[14:11], S_1[14:11], X[14:11], Y[14:11]);
  UBCSuB_17_15 U1 (Co_0, Co_1, So_0, So_1, X[17:15], Y[17:15]);
endmodule

module UBHCSuB_17_4(C, S, X, Y, Ci);
  output C;
  output [17:4] S;
  input Ci;
  input [17:4] X;
  input [17:4] Y;
  wire C_0;
  wire C_1;
  wire Co;
  wire [17:11] S_0;
  wire [17:11] S_1;
  assign S[11] = ( S_0[11] & ( ~ Co ) ) | ( S_1[11] & Co );
  assign S[12] = ( S_0[12] & ( ~ Co ) ) | ( S_1[12] & Co );
  assign S[13] = ( S_0[13] & ( ~ Co ) ) | ( S_1[13] & Co );
  assign S[14] = ( S_0[14] & ( ~ Co ) ) | ( S_1[14] & Co );
  assign S[15] = ( S_0[15] & ( ~ Co ) ) | ( S_1[15] & Co );
  assign S[16] = ( S_0[16] & ( ~ Co ) ) | ( S_1[16] & Co );
  assign S[17] = ( S_0[17] & ( ~ Co ) ) | ( S_1[17] & Co );
  assign C = ( C_0 & ( ~ Co ) ) | ( C_1 & Co );
  UBHCSuB_10_4 U0 (Co, S[10:4], X[10:4], Y[10:4], Ci);
  UBCSuB_17_11 U1 (C_0, C_1, S_0, S_1, X[17:11], Y[17:11]);
endmodule

module UBZero_18_18(O);
  output [18:18] O;
  assign O[18] = 0;
endmodule

module UBOne_18(O);
  output O;
  assign O = 1;
endmodule

module UBFA_18(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSuB_18_18(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_18_18 U0 (Ci_0);
  UBOne_18 U1 (Ci_1);
  UBFA_18 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_18 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBZero_19_19(O);
  output [19:19] O;
  assign O[19] = 0;
endmodule

module UBOne_19(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_19_19(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_19_19 U0 (Ci_0);
  UBOne_19 U1 (Ci_1);
  UBFA_19 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_19 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_19_18(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [19:18] S_0;
  output [19:18] S_1;
  input [19:18] X;
  input [19:18] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire So_0;
  wire So_1;
  assign S_0[19] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[19] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_18_18 U0 (Ci_0, Ci_1, S_0[18], S_1[18], X[18], Y[18]);
  UBCSuB_19_19 U1 (Co_0, Co_1, So_0, So_1, X[19], Y[19]);
endmodule

module UBZero_20_20(O);
  output [20:20] O;
  assign O[20] = 0;
endmodule

module UBOne_20(O);
  output O;
  assign O = 1;
endmodule

module UBFA_20(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSuB_20_20(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_20_20 U0 (Ci_0);
  UBOne_20 U1 (Ci_1);
  UBFA_20 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_20 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBZero_21_21(O);
  output [21:21] O;
  assign O[21] = 0;
endmodule

module UBOne_21(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_21_21(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_21_21 U0 (Ci_0);
  UBOne_21 U1 (Ci_1);
  UBFA_21 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_21 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_21_20(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [21:20] S_0;
  output [21:20] S_1;
  input [21:20] X;
  input [21:20] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire So_0;
  wire So_1;
  assign S_0[21] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[21] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_20_20 U0 (Ci_0, Ci_1, S_0[20], S_1[20], X[20], Y[20]);
  UBCSuB_21_21 U1 (Co_0, Co_1, So_0, So_1, X[21], Y[21]);
endmodule

module UBCSuB_21_18(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [21:18] S_0;
  output [21:18] S_1;
  input [21:18] X;
  input [21:18] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [21:20] So_0;
  wire [21:20] So_1;
  assign S_0[20] = ( So_0[20] & ( ~ Ci_0 ) ) | ( So_1[20] & Ci_0 );
  assign S_0[21] = ( So_0[21] & ( ~ Ci_0 ) ) | ( So_1[21] & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[20] = ( So_0[20] & ( ~ Ci_1 ) ) | ( So_1[20] & Ci_1 );
  assign S_1[21] = ( So_0[21] & ( ~ Ci_1 ) ) | ( So_1[21] & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_19_18 U0 (Ci_0, Ci_1, S_0[19:18], S_1[19:18], X[19:18], Y[19:18]);
  UBCSuB_21_20 U1 (Co_0, Co_1, So_0, So_1, X[21:20], Y[21:20]);
endmodule

module UBZero_22_22(O);
  output [22:22] O;
  assign O[22] = 0;
endmodule

module UBOne_22(O);
  output O;
  assign O = 1;
endmodule

module UBFA_22(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSuB_22_22(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_22_22 U0 (Ci_0);
  UBOne_22 U1 (Ci_1);
  UBFA_22 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_22 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBZero_23_23(O);
  output [23:23] O;
  assign O[23] = 0;
endmodule

module UBOne_23(O);
  output O;
  assign O = 1;
endmodule

module UBFA_23(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSuB_23_23(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_23_23 U0 (Ci_0);
  UBOne_23 U1 (Ci_1);
  UBFA_23 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_23 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_23_22(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [23:22] S_0;
  output [23:22] S_1;
  input [23:22] X;
  input [23:22] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire So_0;
  wire So_1;
  assign S_0[23] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[23] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_22_22 U0 (Ci_0, Ci_1, S_0[22], S_1[22], X[22], Y[22]);
  UBCSuB_23_23 U1 (Co_0, Co_1, So_0, So_1, X[23], Y[23]);
endmodule

module UBZero_24_24(O);
  output [24:24] O;
  assign O[24] = 0;
endmodule

module UBOne_24(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_24_24(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_24_24 U0 (Ci_0);
  UBOne_24 U1 (Ci_1);
  UBFA_24 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_24 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_24_22(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [24:22] S_0;
  output [24:22] S_1;
  input [24:22] X;
  input [24:22] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [24:24] So_0;
  wire [24:24] So_1;
  assign S_0[24] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[24] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_23_22 U0 (Ci_0, Ci_1, S_0[23:22], S_1[23:22], X[23:22], Y[23:22]);
  UBCSuB_24_24 U1 (Co_0, Co_1, So_0, So_1, X[24], Y[24]);
endmodule

module UBCSuB_24_18(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [24:18] S_0;
  output [24:18] S_1;
  input [24:18] X;
  input [24:18] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [24:22] So_0;
  wire [24:22] So_1;
  assign S_0[22] = ( So_0[22] & ( ~ Ci_0 ) ) | ( So_1[22] & Ci_0 );
  assign S_0[23] = ( So_0[23] & ( ~ Ci_0 ) ) | ( So_1[23] & Ci_0 );
  assign S_0[24] = ( So_0[24] & ( ~ Ci_0 ) ) | ( So_1[24] & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[22] = ( So_0[22] & ( ~ Ci_1 ) ) | ( So_1[22] & Ci_1 );
  assign S_1[23] = ( So_0[23] & ( ~ Ci_1 ) ) | ( So_1[23] & Ci_1 );
  assign S_1[24] = ( So_0[24] & ( ~ Ci_1 ) ) | ( So_1[24] & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_21_18 U0 (Ci_0, Ci_1, S_0[21:18], S_1[21:18], X[21:18], Y[21:18]);
  UBCSuB_24_22 U1 (Co_0, Co_1, So_0, So_1, X[24:22], Y[24:22]);
endmodule

module UBZero_25_25(O);
  output [25:25] O;
  assign O[25] = 0;
endmodule

module UBOne_25(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_25_25(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_25_25 U0 (Ci_0);
  UBOne_25 U1 (Ci_1);
  UBFA_25 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_25 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBZero_26_26(O);
  output [26:26] O;
  assign O[26] = 0;
endmodule

module UBOne_26(O);
  output O;
  assign O = 1;
endmodule

module UBFA_26(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSuB_26_26(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_26_26 U0 (Ci_0);
  UBOne_26 U1 (Ci_1);
  UBFA_26 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_26 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_26_25(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [26:25] S_0;
  output [26:25] S_1;
  input [26:25] X;
  input [26:25] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire So_0;
  wire So_1;
  assign S_0[26] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[26] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_25_25 U0 (Ci_0, Ci_1, S_0[25], S_1[25], X[25], Y[25]);
  UBCSuB_26_26 U1 (Co_0, Co_1, So_0, So_1, X[26], Y[26]);
endmodule

module UBZero_27_27(O);
  output [27:27] O;
  assign O[27] = 0;
endmodule

module UBOne_27(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_27_27(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_27_27 U0 (Ci_0);
  UBOne_27 U1 (Ci_1);
  UBFA_27 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_27 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBZero_28_28(O);
  output [28:28] O;
  assign O[28] = 0;
endmodule

module UBOne_28(O);
  output O;
  assign O = 1;
endmodule

module UBFA_28(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSuB_28_28(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_28_28 U0 (Ci_0);
  UBOne_28 U1 (Ci_1);
  UBFA_28 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_28 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_28_27(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [28:27] S_0;
  output [28:27] S_1;
  input [28:27] X;
  input [28:27] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire So_0;
  wire So_1;
  assign S_0[28] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[28] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_27_27 U0 (Ci_0, Ci_1, S_0[27], S_1[27], X[27], Y[27]);
  UBCSuB_28_28 U1 (Co_0, Co_1, So_0, So_1, X[28], Y[28]);
endmodule

module UBCSuB_28_25(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [28:25] S_0;
  output [28:25] S_1;
  input [28:25] X;
  input [28:25] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [28:27] So_0;
  wire [28:27] So_1;
  assign S_0[27] = ( So_0[27] & ( ~ Ci_0 ) ) | ( So_1[27] & Ci_0 );
  assign S_0[28] = ( So_0[28] & ( ~ Ci_0 ) ) | ( So_1[28] & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[27] = ( So_0[27] & ( ~ Ci_1 ) ) | ( So_1[27] & Ci_1 );
  assign S_1[28] = ( So_0[28] & ( ~ Ci_1 ) ) | ( So_1[28] & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_26_25 U0 (Ci_0, Ci_1, S_0[26:25], S_1[26:25], X[26:25], Y[26:25]);
  UBCSuB_28_27 U1 (Co_0, Co_1, So_0, So_1, X[28:27], Y[28:27]);
endmodule

module UBZero_29_29(O);
  output [29:29] O;
  assign O[29] = 0;
endmodule

module UBOne_29(O);
  output O;
  assign O = 1;
endmodule

module UBCSuB_29_29(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_29_29 U0 (Ci_0);
  UBOne_29 U1 (Ci_1);
  UBFA_29 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_29 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBZero_30_30(O);
  output [30:30] O;
  assign O[30] = 0;
endmodule

module UBOne_30(O);
  output O;
  assign O = 1;
endmodule

module UBFA_30(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSuB_30_30(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_30_30 U0 (Ci_0);
  UBOne_30 U1 (Ci_1);
  UBFA_30 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_30 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_30_29(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [30:29] S_0;
  output [30:29] S_1;
  input [30:29] X;
  input [30:29] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire So_0;
  wire So_1;
  assign S_0[30] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[30] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_29_29 U0 (Ci_0, Ci_1, S_0[29], S_1[29], X[29], Y[29]);
  UBCSuB_30_30 U1 (Co_0, Co_1, So_0, So_1, X[30], Y[30]);
endmodule

module UBZero_31_31(O);
  output [31:31] O;
  assign O[31] = 0;
endmodule

module UBOne_31(O);
  output O;
  assign O = 1;
endmodule

module UBFA_31(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSuB_31_31(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output S_0;
  output S_1;
  input X;
  input Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBZero_31_31 U0 (Ci_0);
  UBOne_31 U1 (Ci_1);
  UBFA_31 U2 (Co_0, S_0, X, Y, Ci_0);
  UBFA_31 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBCSuB_31_29(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [31:29] S_0;
  output [31:29] S_1;
  input [31:29] X;
  input [31:29] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [31:31] So_0;
  wire [31:31] So_1;
  assign S_0[31] = ( So_0 & ( ~ Ci_0 ) ) | ( So_1 & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[31] = ( So_0 & ( ~ Ci_1 ) ) | ( So_1 & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_30_29 U0 (Ci_0, Ci_1, S_0[30:29], S_1[30:29], X[30:29], Y[30:29]);
  UBCSuB_31_31 U1 (Co_0, Co_1, So_0, So_1, X[31], Y[31]);
endmodule

module UBCSuB_31_25(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [31:25] S_0;
  output [31:25] S_1;
  input [31:25] X;
  input [31:25] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [31:29] So_0;
  wire [31:29] So_1;
  assign S_0[29] = ( So_0[29] & ( ~ Ci_0 ) ) | ( So_1[29] & Ci_0 );
  assign S_0[30] = ( So_0[30] & ( ~ Ci_0 ) ) | ( So_1[30] & Ci_0 );
  assign S_0[31] = ( So_0[31] & ( ~ Ci_0 ) ) | ( So_1[31] & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[29] = ( So_0[29] & ( ~ Ci_1 ) ) | ( So_1[29] & Ci_1 );
  assign S_1[30] = ( So_0[30] & ( ~ Ci_1 ) ) | ( So_1[30] & Ci_1 );
  assign S_1[31] = ( So_0[31] & ( ~ Ci_1 ) ) | ( So_1[31] & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_28_25 U0 (Ci_0, Ci_1, S_0[28:25], S_1[28:25], X[28:25], Y[28:25]);
  UBCSuB_31_29 U1 (Co_0, Co_1, So_0, So_1, X[31:29], Y[31:29]);
endmodule

module UBCSuB_31_18(C_0, C_1, S_0, S_1, X, Y);
  output C_0;
  output C_1;
  output [31:18] S_0;
  output [31:18] S_1;
  input [31:18] X;
  input [31:18] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [31:25] So_0;
  wire [31:25] So_1;
  assign S_0[25] = ( So_0[25] & ( ~ Ci_0 ) ) | ( So_1[25] & Ci_0 );
  assign S_0[26] = ( So_0[26] & ( ~ Ci_0 ) ) | ( So_1[26] & Ci_0 );
  assign S_0[27] = ( So_0[27] & ( ~ Ci_0 ) ) | ( So_1[27] & Ci_0 );
  assign S_0[28] = ( So_0[28] & ( ~ Ci_0 ) ) | ( So_1[28] & Ci_0 );
  assign S_0[29] = ( So_0[29] & ( ~ Ci_0 ) ) | ( So_1[29] & Ci_0 );
  assign S_0[30] = ( So_0[30] & ( ~ Ci_0 ) ) | ( So_1[30] & Ci_0 );
  assign S_0[31] = ( So_0[31] & ( ~ Ci_0 ) ) | ( So_1[31] & Ci_0 );
  assign C_0 = ( Co_0 & ( ~ Ci_0 ) ) | ( Co_1 & Ci_0 );
  assign S_1[25] = ( So_0[25] & ( ~ Ci_1 ) ) | ( So_1[25] & Ci_1 );
  assign S_1[26] = ( So_0[26] & ( ~ Ci_1 ) ) | ( So_1[26] & Ci_1 );
  assign S_1[27] = ( So_0[27] & ( ~ Ci_1 ) ) | ( So_1[27] & Ci_1 );
  assign S_1[28] = ( So_0[28] & ( ~ Ci_1 ) ) | ( So_1[28] & Ci_1 );
  assign S_1[29] = ( So_0[29] & ( ~ Ci_1 ) ) | ( So_1[29] & Ci_1 );
  assign S_1[30] = ( So_0[30] & ( ~ Ci_1 ) ) | ( So_1[30] & Ci_1 );
  assign S_1[31] = ( So_0[31] & ( ~ Ci_1 ) ) | ( So_1[31] & Ci_1 );
  assign C_1 = ( Co_0 & ( ~ Ci_1 ) ) | ( Co_1 & Ci_1 );
  UBCSuB_24_18 U0 (Ci_0, Ci_1, S_0[24:18], S_1[24:18], X[24:18], Y[24:18]);
  UBCSuB_31_25 U1 (Co_0, Co_1, So_0, So_1, X[31:25], Y[31:25]);
endmodule

module UBPriCSuA_31_4(S, X, Y, Cin);
  output [32:4] S;
  input Cin;
  input [31:4] X;
  input [31:4] Y;
  wire C_0;
  wire C_1;
  wire Co;
  wire [31:18] S_0;
  wire [31:18] S_1;
  assign S[18] = ( S_0[18] & ( ~ Co ) ) | ( S_1[18] & Co );
  assign S[19] = ( S_0[19] & ( ~ Co ) ) | ( S_1[19] & Co );
  assign S[20] = ( S_0[20] & ( ~ Co ) ) | ( S_1[20] & Co );
  assign S[21] = ( S_0[21] & ( ~ Co ) ) | ( S_1[21] & Co );
  assign S[22] = ( S_0[22] & ( ~ Co ) ) | ( S_1[22] & Co );
  assign S[23] = ( S_0[23] & ( ~ Co ) ) | ( S_1[23] & Co );
  assign S[24] = ( S_0[24] & ( ~ Co ) ) | ( S_1[24] & Co );
  assign S[25] = ( S_0[25] & ( ~ Co ) ) | ( S_1[25] & Co );
  assign S[26] = ( S_0[26] & ( ~ Co ) ) | ( S_1[26] & Co );
  assign S[27] = ( S_0[27] & ( ~ Co ) ) | ( S_1[27] & Co );
  assign S[28] = ( S_0[28] & ( ~ Co ) ) | ( S_1[28] & Co );
  assign S[29] = ( S_0[29] & ( ~ Co ) ) | ( S_1[29] & Co );
  assign S[30] = ( S_0[30] & ( ~ Co ) ) | ( S_1[30] & Co );
  assign S[31] = ( S_0[31] & ( ~ Co ) ) | ( S_1[31] & Co );
  assign S[32] = ( C_0 & ( ~ Co ) ) | ( C_1 & Co );
  UBHCSuB_17_4 U0 (Co, S[17:4], X[17:4], Y[17:4], Cin);
  UBCSuB_31_18 U1 (C_0, C_1, S_0, S_1, X[31:18], Y[31:18]);
endmodule

module UBZero_4_4(O);
  output [4:4] O;
  assign O[4] = 0;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module Multiplier_15_0_1000(P, IN1, IN2);
  output [31:0] P;
  input [15:0] IN1;
  input [15:0] IN2;
  wire [32:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  assign P[12] = W[12];
  assign P[13] = W[13];
  assign P[14] = W[14];
  assign P[15] = W[15];
  assign P[16] = W[16];
  assign P[17] = W[17];
  assign P[18] = W[18];
  assign P[19] = W[19];
  assign P[20] = W[20];
  assign P[21] = W[21];
  assign P[22] = W[22];
  assign P[23] = W[23];
  assign P[24] = W[24];
  assign P[25] = W[25];
  assign P[26] = W[26];
  assign P[27] = W[27];
  assign P[28] = W[28];
  assign P[29] = W[29];
  assign P[30] = W[30];
  assign P[31] = W[31];
  MultUB_STD_C42_CS000 U0 (W, IN1, IN2);
endmodule

module C42TR_15_0_16_1_1000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15);
  output [31:4] S1;
  output [31:0] S2;
  input [15:0] PP0;
  input [16:1] PP1;
  input [25:10] PP10;
  input [26:11] PP11;
  input [27:12] PP12;
  input [28:13] PP13;
  input [29:14] PP14;
  input [30:15] PP15;
  input [17:2] PP2;
  input [18:3] PP3;
  input [19:4] PP4;
  input [20:5] PP5;
  input [21:6] PP6;
  input [22:7] PP7;
  input [23:8] PP8;
  input [24:9] PP9;
  wire [18:0] W1_0;
  wire [18:2] W1_1;
  wire [22:4] W1_2;
  wire [22:6] W1_3;
  wire [26:8] W1_4;
  wire [26:10] W1_5;
  wire [30:12] W1_6;
  wire [30:14] W1_7;
  wire [30:8] W2_10;
  wire [31:11] W2_11;
  wire [22:0] W2_8;
  wire [23:3] W2_9;
  UB4_2Comp_15_0_16000 U0 (W1_1[18:2], W1_0[18:0], PP0, PP1, PP2, PP3);
  UB4_2Comp_19_4_20000 U1 (W1_3[22:6], W1_2[22:4], PP4, PP5, PP6, PP7);
  UB4_2Comp_23_8_24000 U2 (W1_5[26:10], W1_4[26:8], PP8, PP9, PP10, PP11);
  UB4_2Comp_27_12_2000 U3 (W1_7[30:14], W1_6[30:12], PP12, PP13, PP14, PP15);
  UB4_2Comp_18_0_18000 U4 (W2_9[23:3], W2_8[22:0], W1_0[18:0], W1_1[18:2], W1_2[22:4], W1_3[22:6]);
  UB4_2Comp_26_8_26000 U5 (W2_11[31:11], W2_10[30:8], W1_4[26:8], W1_5[26:10], W1_6[30:12], W1_7[30:14]);
  UB4_2Comp_22_0_23000 U6 (S1[31:4], S2[31:0], W2_8[22:0], W2_9[23:3], W2_10[30:8], W2_11[31:11]);
endmodule

module MultUB_STD_C42_CS000 (P, IN1, IN2);
  output [32:0] P;
  input [15:0] IN1;
  input [15:0] IN2;
  wire [15:0] PP0;
  wire [16:1] PP1;
  wire [25:10] PP10;
  wire [26:11] PP11;
  wire [27:12] PP12;
  wire [28:13] PP13;
  wire [29:14] PP14;
  wire [30:15] PP15;
  wire [17:2] PP2;
  wire [18:3] PP3;
  wire [19:4] PP4;
  wire [20:5] PP5;
  wire [21:6] PP6;
  wire [22:7] PP7;
  wire [23:8] PP8;
  wire [24:9] PP9;
  wire [31:4] S1;
  wire [31:0] S2;
  UBPPG_15_0_15_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, IN1, IN2);
  C42TR_15_0_16_1_1000 U1 (S1[31:4], S2[31:0], PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15);
  UBCSu_31_4_31_0 U2 (P, S1[31:4], S2[31:0]);
endmodule

module PureCSA_10_8 (C, S, X, Y, Z);
  output [11:9] C;
  output [10:8] S;
  input [10:8] X;
  input [10:8] Y;
  input [10:8] Z;
  UBFA_8 U0 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U1 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U2 (C[11], S[10], X[10], Y[10], Z[10]);
endmodule

module PureCSA_13_12 (C, S, X, Y, Z);
  output [14:13] C;
  output [13:12] S;
  input [13:12] X;
  input [13:12] Y;
  input [13:12] Z;
  UBFA_12 U0 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U1 (C[14], S[13], X[13], Y[13], Z[13]);
endmodule

module PureCSA_5_4 (C, S, X, Y, Z);
  output [6:5] C;
  output [5:4] S;
  input [5:4] X;
  input [5:4] Y;
  input [5:4] Z;
  UBFA_4 U0 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U1 (C[6], S[5], X[5], Y[5], Z[5]);
endmodule

module PureCSHA_11_10 (C, S, X, Y);
  output [12:11] C;
  output [11:10] S;
  input [11:10] X;
  input [11:10] Y;
  UBHA_10 U0 (C[11], S[10], X[10], Y[10]);
  UBHA_11 U1 (C[12], S[11], X[11], Y[11]);
endmodule

module PureCSHA_22_20 (C, S, X, Y);
  output [23:21] C;
  output [22:20] S;
  input [22:20] X;
  input [22:20] Y;
  UBHA_20 U0 (C[21], S[20], X[20], Y[20]);
  UBHA_21 U1 (C[22], S[21], X[21], Y[21]);
  UBHA_22 U2 (C[23], S[22], X[22], Y[22]);
endmodule

module PureCSHA_30_25 (C, S, X, Y);
  output [31:26] C;
  output [30:25] S;
  input [30:25] X;
  input [30:25] Y;
  UBHA_25 U0 (C[26], S[25], X[25], Y[25]);
  UBHA_26 U1 (C[27], S[26], X[26], Y[26]);
  UBHA_27 U2 (C[28], S[27], X[27], Y[27]);
  UBHA_28 U3 (C[29], S[28], X[28], Y[28]);
  UBHA_29 U4 (C[30], S[29], X[29], Y[29]);
  UBHA_30 U5 (C[31], S[30], X[30], Y[30]);
endmodule

module PureCSHA_30_28 (C, S, X, Y);
  output [31:29] C;
  output [30:28] S;
  input [30:28] X;
  input [30:28] Y;
  UBHA_28 U0 (C[29], S[28], X[28], Y[28]);
  UBHA_29 U1 (C[30], S[29], X[29], Y[29]);
  UBHA_30 U2 (C[31], S[30], X[30], Y[30]);
endmodule

module PureCSHA_3_2 (C, S, X, Y);
  output [4:3] C;
  output [3:2] S;
  input [3:2] X;
  input [3:2] Y;
  UBHA_2 U0 (C[3], S[2], X[2], Y[2]);
  UBHA_3 U1 (C[4], S[3], X[3], Y[3]);
endmodule

module PureCSHA_7_3 (C, S, X, Y);
  output [8:4] C;
  output [7:3] S;
  input [7:3] X;
  input [7:3] Y;
  UBHA_3 U0 (C[4], S[3], X[3], Y[3]);
  UBHA_4 U1 (C[5], S[4], X[4], Y[4]);
  UBHA_5 U2 (C[6], S[5], X[5], Y[5]);
  UBHA_6 U3 (C[7], S[6], X[6], Y[6]);
  UBHA_7 U4 (C[8], S[7], X[7], Y[7]);
endmodule

module UB4_2Comp_15_0_16000 (C, S, IN0, IN1, IN2, IN3);
  output [18:2] C;
  output [18:0] S;
  input [15:0] IN0;
  input [16:1] IN1;
  input [17:2] IN2;
  input [18:3] IN3;
  wire W0;
  wire W1;
  wire WZ;
  UB1DCON_0 U0 (S[0], IN0[0]);
  UBHA_1 U1 (C[2], S[1], IN1[1], IN0[1]);
  UBFA_2 U2 (C[3], S[2], IN2[2], IN1[2], IN0[2]);
  UBZero_3_3 U3 (WZ);
  UBPure4_2CMP_15_3 U4 (W0, C[16:4], S[15:3], IN3[15:3], IN2[15:3], IN1[15:3], IN0[15:3], WZ);
  UB1B3_2CMP_16 U5 (W1, C[17], S[16], IN3[16], IN2[16], IN1[16], W0);
  UBFA_17 U6 (C[18], S[17], IN3[17], IN2[17], W1);
  UB1DCON_18 U7 (S[18], IN3[18]);
endmodule

module UB4_2Comp_18_0_18000 (C, S, IN0, IN1, IN2, IN3);
  output [23:3] C;
  output [22:0] S;
  input [18:0] IN0;
  input [18:2] IN1;
  input [22:4] IN2;
  input [22:6] IN3;
  wire W0;
  wire WZ;
  UBCON_1_0 U0 (S[1:0], IN0[1:0]);
  PureCSHA_3_2 U1 (C[4:3], S[3:2], IN1[3:2], IN0[3:2]);
  PureCSA_5_4 U2 (C[6:5], S[5:4], IN2[5:4], IN1[5:4], IN0[5:4]);
  UBZero_6_6 U3 (WZ);
  UBPure4_2CMP_18_6 U4 (W0, C[19:7], S[18:6], IN3[18:6], IN2[18:6], IN1[18:6], IN0[18:6], WZ);
  UBFA_19 U5 (C[20], S[19], IN3[19], IN2[19], W0);
  PureCSHA_22_20 U6 (C[23:21], S[22:20], IN3[22:20], IN2[22:20]);
endmodule

module UB4_2Comp_19_4_20000 (C, S, IN0, IN1, IN2, IN3);
  output [22:6] C;
  output [22:4] S;
  input [19:4] IN0;
  input [20:5] IN1;
  input [21:6] IN2;
  input [22:7] IN3;
  wire W0;
  wire W1;
  wire WZ;
  UB1DCON_4 U0 (S[4], IN0[4]);
  UBHA_5 U1 (C[6], S[5], IN1[5], IN0[5]);
  UBFA_6 U2 (C[7], S[6], IN2[6], IN1[6], IN0[6]);
  UBZero_7_7 U3 (WZ);
  UBPure4_2CMP_19_7 U4 (W0, C[20:8], S[19:7], IN3[19:7], IN2[19:7], IN1[19:7], IN0[19:7], WZ);
  UB1B3_2CMP_20 U5 (W1, C[21], S[20], IN3[20], IN2[20], IN1[20], W0);
  UBFA_21 U6 (C[22], S[21], IN3[21], IN2[21], W1);
  UB1DCON_22 U7 (S[22], IN3[22]);
endmodule

module UB4_2Comp_22_0_23000 (C, S, IN0, IN1, IN2, IN3);
  output [31:4] C;
  output [31:0] S;
  input [22:0] IN0;
  input [23:3] IN1;
  input [30:8] IN2;
  input [31:11] IN3;
  wire W0;
  wire W1;
  wire WZ;
  UBCON_2_0 U0 (S[2:0], IN0[2:0]);
  PureCSHA_7_3 U1 (C[8:4], S[7:3], IN1[7:3], IN0[7:3]);
  PureCSA_10_8 U2 (C[11:9], S[10:8], IN2[10:8], IN1[10:8], IN0[10:8]);
  UBZero_11_11 U3 (WZ);
  UBPure4_2CMP_22_1000 U4 (W0, C[23:12], S[22:11], IN3[22:11], IN2[22:11], IN1[22:11], IN0[22:11], WZ);
  UB1B3_2CMP_23 U5 (W1, C[24], S[23], IN3[23], IN2[23], IN1[23], W0);
  UBFA_24 U6 (C[25], S[24], IN3[24], IN2[24], W1);
  PureCSHA_30_25 U7 (C[31:26], S[30:25], IN3[30:25], IN2[30:25]);
  UB1DCON_31 U8 (S[31], IN3[31]);
endmodule

module UB4_2Comp_23_8_24000 (C, S, IN0, IN1, IN2, IN3);
  output [26:10] C;
  output [26:8] S;
  input [23:8] IN0;
  input [24:9] IN1;
  input [25:10] IN2;
  input [26:11] IN3;
  wire W0;
  wire W1;
  wire WZ;
  UB1DCON_8 U0 (S[8], IN0[8]);
  UBHA_9 U1 (C[10], S[9], IN1[9], IN0[9]);
  UBFA_10 U2 (C[11], S[10], IN2[10], IN1[10], IN0[10]);
  UBZero_11_11 U3 (WZ);
  UBPure4_2CMP_23_1000 U4 (W0, C[24:12], S[23:11], IN3[23:11], IN2[23:11], IN1[23:11], IN0[23:11], WZ);
  UB1B3_2CMP_24 U5 (W1, C[25], S[24], IN3[24], IN2[24], IN1[24], W0);
  UBFA_25 U6 (C[26], S[25], IN3[25], IN2[25], W1);
  UB1DCON_26 U7 (S[26], IN3[26]);
endmodule

module UB4_2Comp_26_8_26000 (C, S, IN0, IN1, IN2, IN3);
  output [31:11] C;
  output [30:8] S;
  input [26:8] IN0;
  input [26:10] IN1;
  input [30:12] IN2;
  input [30:14] IN3;
  wire W0;
  wire WZ;
  UBCON_9_8 U0 (S[9:8], IN0[9:8]);
  PureCSHA_11_10 U1 (C[12:11], S[11:10], IN1[11:10], IN0[11:10]);
  PureCSA_13_12 U2 (C[14:13], S[13:12], IN2[13:12], IN1[13:12], IN0[13:12]);
  UBZero_14_14 U3 (WZ);
  UBPure4_2CMP_26_1000 U4 (W0, C[27:15], S[26:14], IN3[26:14], IN2[26:14], IN1[26:14], IN0[26:14], WZ);
  UBFA_27 U5 (C[28], S[27], IN3[27], IN2[27], W0);
  PureCSHA_30_28 U6 (C[31:29], S[30:28], IN3[30:28], IN2[30:28]);
endmodule

module UB4_2Comp_27_12_2000 (C, S, IN0, IN1, IN2, IN3);
  output [30:14] C;
  output [30:12] S;
  input [27:12] IN0;
  input [28:13] IN1;
  input [29:14] IN2;
  input [30:15] IN3;
  wire W0;
  wire W1;
  wire WZ;
  UB1DCON_12 U0 (S[12], IN0[12]);
  UBHA_13 U1 (C[14], S[13], IN1[13], IN0[13]);
  UBFA_14 U2 (C[15], S[14], IN2[14], IN1[14], IN0[14]);
  UBZero_15_15 U3 (WZ);
  UBPure4_2CMP_27_1000 U4 (W0, C[28:16], S[27:15], IN3[27:15], IN2[27:15], IN1[27:15], IN0[27:15], WZ);
  UB1B3_2CMP_28 U5 (W1, C[29], S[28], IN3[28], IN2[28], IN1[28], W0);
  UBFA_29 U6 (C[30], S[29], IN3[29], IN2[29], W1);
  UB1DCON_30 U7 (S[30], IN3[30]);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBCON_3_0 (O, I);
  output [3:0] O;
  input [3:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
endmodule

module UBCON_9_8 (O, I);
  output [9:8] O;
  input [9:8] I;
  UB1DCON_8 U0 (O[8], I[8]);
  UB1DCON_9 U1 (O[9], I[9]);
endmodule

module UBCSu_31_4_31_0 (S, X, Y);
  output [32:0] S;
  input [31:4] X;
  input [31:0] Y;
  UBPureCSu_31_4 U0 (S[32:4], X[31:4], Y[31:4]);
  UBCON_3_0 U1 (S[3:0], Y[3:0]);
endmodule

module UBPPG_15_0_15_0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, IN1, IN2);
  output [15:0] PP0;
  output [16:1] PP1;
  output [25:10] PP10;
  output [26:11] PP11;
  output [27:12] PP12;
  output [28:13] PP13;
  output [29:14] PP14;
  output [30:15] PP15;
  output [17:2] PP2;
  output [18:3] PP3;
  output [19:4] PP4;
  output [20:5] PP5;
  output [21:6] PP6;
  output [22:7] PP7;
  output [23:8] PP8;
  output [24:9] PP9;
  input [15:0] IN1;
  input [15:0] IN2;
  UBVPPG_15_0_0 U0 (PP0, IN1, IN2[0]);
  UBVPPG_15_0_1 U1 (PP1, IN1, IN2[1]);
  UBVPPG_15_0_2 U2 (PP2, IN1, IN2[2]);
  UBVPPG_15_0_3 U3 (PP3, IN1, IN2[3]);
  UBVPPG_15_0_4 U4 (PP4, IN1, IN2[4]);
  UBVPPG_15_0_5 U5 (PP5, IN1, IN2[5]);
  UBVPPG_15_0_6 U6 (PP6, IN1, IN2[6]);
  UBVPPG_15_0_7 U7 (PP7, IN1, IN2[7]);
  UBVPPG_15_0_8 U8 (PP8, IN1, IN2[8]);
  UBVPPG_15_0_9 U9 (PP9, IN1, IN2[9]);
  UBVPPG_15_0_10 U10 (PP10, IN1, IN2[10]);
  UBVPPG_15_0_11 U11 (PP11, IN1, IN2[11]);
  UBVPPG_15_0_12 U12 (PP12, IN1, IN2[12]);
  UBVPPG_15_0_13 U13 (PP13, IN1, IN2[13]);
  UBVPPG_15_0_14 U14 (PP14, IN1, IN2[14]);
  UBVPPG_15_0_15 U15 (PP15, IN1, IN2[15]);
endmodule

module UBPure4_2CMP_15_3 (Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output [16:4] C;
  output Co;
  output [15:3] S;
  input Ci;
  input [15:3] IN0;
  input [15:3] IN1;
  input [15:3] IN2;
  input [15:3] IN3;
  wire [15:4] W;
  UB1B4_2CMP_3 U0 (W[4], C[4], S[3], IN0[3], IN1[3], IN2[3], IN3[3], Ci);
  UB1B4_2CMP_4 U1 (W[5], C[5], S[4], IN0[4], IN1[4], IN2[4], IN3[4], W[4]);
  UB1B4_2CMP_5 U2 (W[6], C[6], S[5], IN0[5], IN1[5], IN2[5], IN3[5], W[5]);
  UB1B4_2CMP_6 U3 (W[7], C[7], S[6], IN0[6], IN1[6], IN2[6], IN3[6], W[6]);
  UB1B4_2CMP_7 U4 (W[8], C[8], S[7], IN0[7], IN1[7], IN2[7], IN3[7], W[7]);
  UB1B4_2CMP_8 U5 (W[9], C[9], S[8], IN0[8], IN1[8], IN2[8], IN3[8], W[8]);
  UB1B4_2CMP_9 U6 (W[10], C[10], S[9], IN0[9], IN1[9], IN2[9], IN3[9], W[9]);
  UB1B4_2CMP_10 U7 (W[11], C[11], S[10], IN0[10], IN1[10], IN2[10], IN3[10], W[10]);
  UB1B4_2CMP_11 U8 (W[12], C[12], S[11], IN0[11], IN1[11], IN2[11], IN3[11], W[11]);
  UB1B4_2CMP_12 U9 (W[13], C[13], S[12], IN0[12], IN1[12], IN2[12], IN3[12], W[12]);
  UB1B4_2CMP_13 U10 (W[14], C[14], S[13], IN0[13], IN1[13], IN2[13], IN3[13], W[13]);
  UB1B4_2CMP_14 U11 (W[15], C[15], S[14], IN0[14], IN1[14], IN2[14], IN3[14], W[14]);
  UB1B4_2CMP_15 U12 (Co, C[16], S[15], IN0[15], IN1[15], IN2[15], IN3[15], W[15]);
endmodule

module UBPure4_2CMP_18_6 (Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output [19:7] C;
  output Co;
  output [18:6] S;
  input Ci;
  input [18:6] IN0;
  input [18:6] IN1;
  input [18:6] IN2;
  input [18:6] IN3;
  wire [18:7] W;
  UB1B4_2CMP_6 U0 (W[7], C[7], S[6], IN0[6], IN1[6], IN2[6], IN3[6], Ci);
  UB1B4_2CMP_7 U1 (W[8], C[8], S[7], IN0[7], IN1[7], IN2[7], IN3[7], W[7]);
  UB1B4_2CMP_8 U2 (W[9], C[9], S[8], IN0[8], IN1[8], IN2[8], IN3[8], W[8]);
  UB1B4_2CMP_9 U3 (W[10], C[10], S[9], IN0[9], IN1[9], IN2[9], IN3[9], W[9]);
  UB1B4_2CMP_10 U4 (W[11], C[11], S[10], IN0[10], IN1[10], IN2[10], IN3[10], W[10]);
  UB1B4_2CMP_11 U5 (W[12], C[12], S[11], IN0[11], IN1[11], IN2[11], IN3[11], W[11]);
  UB1B4_2CMP_12 U6 (W[13], C[13], S[12], IN0[12], IN1[12], IN2[12], IN3[12], W[12]);
  UB1B4_2CMP_13 U7 (W[14], C[14], S[13], IN0[13], IN1[13], IN2[13], IN3[13], W[13]);
  UB1B4_2CMP_14 U8 (W[15], C[15], S[14], IN0[14], IN1[14], IN2[14], IN3[14], W[14]);
  UB1B4_2CMP_15 U9 (W[16], C[16], S[15], IN0[15], IN1[15], IN2[15], IN3[15], W[15]);
  UB1B4_2CMP_16 U10 (W[17], C[17], S[16], IN0[16], IN1[16], IN2[16], IN3[16], W[16]);
  UB1B4_2CMP_17 U11 (W[18], C[18], S[17], IN0[17], IN1[17], IN2[17], IN3[17], W[17]);
  UB1B4_2CMP_18 U12 (Co, C[19], S[18], IN0[18], IN1[18], IN2[18], IN3[18], W[18]);
endmodule

module UBPure4_2CMP_19_7 (Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output [20:8] C;
  output Co;
  output [19:7] S;
  input Ci;
  input [19:7] IN0;
  input [19:7] IN1;
  input [19:7] IN2;
  input [19:7] IN3;
  wire [19:8] W;
  UB1B4_2CMP_7 U0 (W[8], C[8], S[7], IN0[7], IN1[7], IN2[7], IN3[7], Ci);
  UB1B4_2CMP_8 U1 (W[9], C[9], S[8], IN0[8], IN1[8], IN2[8], IN3[8], W[8]);
  UB1B4_2CMP_9 U2 (W[10], C[10], S[9], IN0[9], IN1[9], IN2[9], IN3[9], W[9]);
  UB1B4_2CMP_10 U3 (W[11], C[11], S[10], IN0[10], IN1[10], IN2[10], IN3[10], W[10]);
  UB1B4_2CMP_11 U4 (W[12], C[12], S[11], IN0[11], IN1[11], IN2[11], IN3[11], W[11]);
  UB1B4_2CMP_12 U5 (W[13], C[13], S[12], IN0[12], IN1[12], IN2[12], IN3[12], W[12]);
  UB1B4_2CMP_13 U6 (W[14], C[14], S[13], IN0[13], IN1[13], IN2[13], IN3[13], W[13]);
  UB1B4_2CMP_14 U7 (W[15], C[15], S[14], IN0[14], IN1[14], IN2[14], IN3[14], W[14]);
  UB1B4_2CMP_15 U8 (W[16], C[16], S[15], IN0[15], IN1[15], IN2[15], IN3[15], W[15]);
  UB1B4_2CMP_16 U9 (W[17], C[17], S[16], IN0[16], IN1[16], IN2[16], IN3[16], W[16]);
  UB1B4_2CMP_17 U10 (W[18], C[18], S[17], IN0[17], IN1[17], IN2[17], IN3[17], W[17]);
  UB1B4_2CMP_18 U11 (W[19], C[19], S[18], IN0[18], IN1[18], IN2[18], IN3[18], W[18]);
  UB1B4_2CMP_19 U12 (Co, C[20], S[19], IN0[19], IN1[19], IN2[19], IN3[19], W[19]);
endmodule

module UBPure4_2CMP_22_1000 (Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output [23:12] C;
  output Co;
  output [22:11] S;
  input Ci;
  input [22:11] IN0;
  input [22:11] IN1;
  input [22:11] IN2;
  input [22:11] IN3;
  wire [22:12] W;
  UB1B4_2CMP_11 U0 (W[12], C[12], S[11], IN0[11], IN1[11], IN2[11], IN3[11], Ci);
  UB1B4_2CMP_12 U1 (W[13], C[13], S[12], IN0[12], IN1[12], IN2[12], IN3[12], W[12]);
  UB1B4_2CMP_13 U2 (W[14], C[14], S[13], IN0[13], IN1[13], IN2[13], IN3[13], W[13]);
  UB1B4_2CMP_14 U3 (W[15], C[15], S[14], IN0[14], IN1[14], IN2[14], IN3[14], W[14]);
  UB1B4_2CMP_15 U4 (W[16], C[16], S[15], IN0[15], IN1[15], IN2[15], IN3[15], W[15]);
  UB1B4_2CMP_16 U5 (W[17], C[17], S[16], IN0[16], IN1[16], IN2[16], IN3[16], W[16]);
  UB1B4_2CMP_17 U6 (W[18], C[18], S[17], IN0[17], IN1[17], IN2[17], IN3[17], W[17]);
  UB1B4_2CMP_18 U7 (W[19], C[19], S[18], IN0[18], IN1[18], IN2[18], IN3[18], W[18]);
  UB1B4_2CMP_19 U8 (W[20], C[20], S[19], IN0[19], IN1[19], IN2[19], IN3[19], W[19]);
  UB1B4_2CMP_20 U9 (W[21], C[21], S[20], IN0[20], IN1[20], IN2[20], IN3[20], W[20]);
  UB1B4_2CMP_21 U10 (W[22], C[22], S[21], IN0[21], IN1[21], IN2[21], IN3[21], W[21]);
  UB1B4_2CMP_22 U11 (Co, C[23], S[22], IN0[22], IN1[22], IN2[22], IN3[22], W[22]);
endmodule

module UBPure4_2CMP_23_1000 (Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output [24:12] C;
  output Co;
  output [23:11] S;
  input Ci;
  input [23:11] IN0;
  input [23:11] IN1;
  input [23:11] IN2;
  input [23:11] IN3;
  wire [23:12] W;
  UB1B4_2CMP_11 U0 (W[12], C[12], S[11], IN0[11], IN1[11], IN2[11], IN3[11], Ci);
  UB1B4_2CMP_12 U1 (W[13], C[13], S[12], IN0[12], IN1[12], IN2[12], IN3[12], W[12]);
  UB1B4_2CMP_13 U2 (W[14], C[14], S[13], IN0[13], IN1[13], IN2[13], IN3[13], W[13]);
  UB1B4_2CMP_14 U3 (W[15], C[15], S[14], IN0[14], IN1[14], IN2[14], IN3[14], W[14]);
  UB1B4_2CMP_15 U4 (W[16], C[16], S[15], IN0[15], IN1[15], IN2[15], IN3[15], W[15]);
  UB1B4_2CMP_16 U5 (W[17], C[17], S[16], IN0[16], IN1[16], IN2[16], IN3[16], W[16]);
  UB1B4_2CMP_17 U6 (W[18], C[18], S[17], IN0[17], IN1[17], IN2[17], IN3[17], W[17]);
  UB1B4_2CMP_18 U7 (W[19], C[19], S[18], IN0[18], IN1[18], IN2[18], IN3[18], W[18]);
  UB1B4_2CMP_19 U8 (W[20], C[20], S[19], IN0[19], IN1[19], IN2[19], IN3[19], W[19]);
  UB1B4_2CMP_20 U9 (W[21], C[21], S[20], IN0[20], IN1[20], IN2[20], IN3[20], W[20]);
  UB1B4_2CMP_21 U10 (W[22], C[22], S[21], IN0[21], IN1[21], IN2[21], IN3[21], W[21]);
  UB1B4_2CMP_22 U11 (W[23], C[23], S[22], IN0[22], IN1[22], IN2[22], IN3[22], W[22]);
  UB1B4_2CMP_23 U12 (Co, C[24], S[23], IN0[23], IN1[23], IN2[23], IN3[23], W[23]);
endmodule

module UBPure4_2CMP_26_1000 (Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output [27:15] C;
  output Co;
  output [26:14] S;
  input Ci;
  input [26:14] IN0;
  input [26:14] IN1;
  input [26:14] IN2;
  input [26:14] IN3;
  wire [26:15] W;
  UB1B4_2CMP_14 U0 (W[15], C[15], S[14], IN0[14], IN1[14], IN2[14], IN3[14], Ci);
  UB1B4_2CMP_15 U1 (W[16], C[16], S[15], IN0[15], IN1[15], IN2[15], IN3[15], W[15]);
  UB1B4_2CMP_16 U2 (W[17], C[17], S[16], IN0[16], IN1[16], IN2[16], IN3[16], W[16]);
  UB1B4_2CMP_17 U3 (W[18], C[18], S[17], IN0[17], IN1[17], IN2[17], IN3[17], W[17]);
  UB1B4_2CMP_18 U4 (W[19], C[19], S[18], IN0[18], IN1[18], IN2[18], IN3[18], W[18]);
  UB1B4_2CMP_19 U5 (W[20], C[20], S[19], IN0[19], IN1[19], IN2[19], IN3[19], W[19]);
  UB1B4_2CMP_20 U6 (W[21], C[21], S[20], IN0[20], IN1[20], IN2[20], IN3[20], W[20]);
  UB1B4_2CMP_21 U7 (W[22], C[22], S[21], IN0[21], IN1[21], IN2[21], IN3[21], W[21]);
  UB1B4_2CMP_22 U8 (W[23], C[23], S[22], IN0[22], IN1[22], IN2[22], IN3[22], W[22]);
  UB1B4_2CMP_23 U9 (W[24], C[24], S[23], IN0[23], IN1[23], IN2[23], IN3[23], W[23]);
  UB1B4_2CMP_24 U10 (W[25], C[25], S[24], IN0[24], IN1[24], IN2[24], IN3[24], W[24]);
  UB1B4_2CMP_25 U11 (W[26], C[26], S[25], IN0[25], IN1[25], IN2[25], IN3[25], W[25]);
  UB1B4_2CMP_26 U12 (Co, C[27], S[26], IN0[26], IN1[26], IN2[26], IN3[26], W[26]);
endmodule

module UBPure4_2CMP_27_1000 (Co, C, S, IN0, IN1, IN2, IN3, Ci);
  output [28:16] C;
  output Co;
  output [27:15] S;
  input Ci;
  input [27:15] IN0;
  input [27:15] IN1;
  input [27:15] IN2;
  input [27:15] IN3;
  wire [27:16] W;
  UB1B4_2CMP_15 U0 (W[16], C[16], S[15], IN0[15], IN1[15], IN2[15], IN3[15], Ci);
  UB1B4_2CMP_16 U1 (W[17], C[17], S[16], IN0[16], IN1[16], IN2[16], IN3[16], W[16]);
  UB1B4_2CMP_17 U2 (W[18], C[18], S[17], IN0[17], IN1[17], IN2[17], IN3[17], W[17]);
  UB1B4_2CMP_18 U3 (W[19], C[19], S[18], IN0[18], IN1[18], IN2[18], IN3[18], W[18]);
  UB1B4_2CMP_19 U4 (W[20], C[20], S[19], IN0[19], IN1[19], IN2[19], IN3[19], W[19]);
  UB1B4_2CMP_20 U5 (W[21], C[21], S[20], IN0[20], IN1[20], IN2[20], IN3[20], W[20]);
  UB1B4_2CMP_21 U6 (W[22], C[22], S[21], IN0[21], IN1[21], IN2[21], IN3[21], W[21]);
  UB1B4_2CMP_22 U7 (W[23], C[23], S[22], IN0[22], IN1[22], IN2[22], IN3[22], W[22]);
  UB1B4_2CMP_23 U8 (W[24], C[24], S[23], IN0[23], IN1[23], IN2[23], IN3[23], W[23]);
  UB1B4_2CMP_24 U9 (W[25], C[25], S[24], IN0[24], IN1[24], IN2[24], IN3[24], W[24]);
  UB1B4_2CMP_25 U10 (W[26], C[26], S[25], IN0[25], IN1[25], IN2[25], IN3[25], W[25]);
  UB1B4_2CMP_26 U11 (W[27], C[27], S[26], IN0[26], IN1[26], IN2[26], IN3[26], W[26]);
  UB1B4_2CMP_27 U12 (Co, C[28], S[27], IN0[27], IN1[27], IN2[27], IN3[27], W[27]);
endmodule

module UBPureCSu_31_4 (S, X, Y);
  output [32:4] S;
  input [31:4] X;
  input [31:4] Y;
  wire C;
  UBPriCSuA_31_4 U0 (S, X, Y, C);
  UBZero_4_4 U1 (C);
endmodule

module UBVPPG_15_0_0 (O, IN1, IN2);
  output [15:0] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
  UB1BPPG_6_0 U6 (O[6], IN1[6], IN2);
  UB1BPPG_7_0 U7 (O[7], IN1[7], IN2);
  UB1BPPG_8_0 U8 (O[8], IN1[8], IN2);
  UB1BPPG_9_0 U9 (O[9], IN1[9], IN2);
  UB1BPPG_10_0 U10 (O[10], IN1[10], IN2);
  UB1BPPG_11_0 U11 (O[11], IN1[11], IN2);
  UB1BPPG_12_0 U12 (O[12], IN1[12], IN2);
  UB1BPPG_13_0 U13 (O[13], IN1[13], IN2);
  UB1BPPG_14_0 U14 (O[14], IN1[14], IN2);
  UB1BPPG_15_0 U15 (O[15], IN1[15], IN2);
endmodule

module UBVPPG_15_0_1 (O, IN1, IN2);
  output [16:1] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_1 U0 (O[1], IN1[0], IN2);
  UB1BPPG_1_1 U1 (O[2], IN1[1], IN2);
  UB1BPPG_2_1 U2 (O[3], IN1[2], IN2);
  UB1BPPG_3_1 U3 (O[4], IN1[3], IN2);
  UB1BPPG_4_1 U4 (O[5], IN1[4], IN2);
  UB1BPPG_5_1 U5 (O[6], IN1[5], IN2);
  UB1BPPG_6_1 U6 (O[7], IN1[6], IN2);
  UB1BPPG_7_1 U7 (O[8], IN1[7], IN2);
  UB1BPPG_8_1 U8 (O[9], IN1[8], IN2);
  UB1BPPG_9_1 U9 (O[10], IN1[9], IN2);
  UB1BPPG_10_1 U10 (O[11], IN1[10], IN2);
  UB1BPPG_11_1 U11 (O[12], IN1[11], IN2);
  UB1BPPG_12_1 U12 (O[13], IN1[12], IN2);
  UB1BPPG_13_1 U13 (O[14], IN1[13], IN2);
  UB1BPPG_14_1 U14 (O[15], IN1[14], IN2);
  UB1BPPG_15_1 U15 (O[16], IN1[15], IN2);
endmodule

module UBVPPG_15_0_10 (O, IN1, IN2);
  output [25:10] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_10 U0 (O[10], IN1[0], IN2);
  UB1BPPG_1_10 U1 (O[11], IN1[1], IN2);
  UB1BPPG_2_10 U2 (O[12], IN1[2], IN2);
  UB1BPPG_3_10 U3 (O[13], IN1[3], IN2);
  UB1BPPG_4_10 U4 (O[14], IN1[4], IN2);
  UB1BPPG_5_10 U5 (O[15], IN1[5], IN2);
  UB1BPPG_6_10 U6 (O[16], IN1[6], IN2);
  UB1BPPG_7_10 U7 (O[17], IN1[7], IN2);
  UB1BPPG_8_10 U8 (O[18], IN1[8], IN2);
  UB1BPPG_9_10 U9 (O[19], IN1[9], IN2);
  UB1BPPG_10_10 U10 (O[20], IN1[10], IN2);
  UB1BPPG_11_10 U11 (O[21], IN1[11], IN2);
  UB1BPPG_12_10 U12 (O[22], IN1[12], IN2);
  UB1BPPG_13_10 U13 (O[23], IN1[13], IN2);
  UB1BPPG_14_10 U14 (O[24], IN1[14], IN2);
  UB1BPPG_15_10 U15 (O[25], IN1[15], IN2);
endmodule

module UBVPPG_15_0_11 (O, IN1, IN2);
  output [26:11] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_11 U0 (O[11], IN1[0], IN2);
  UB1BPPG_1_11 U1 (O[12], IN1[1], IN2);
  UB1BPPG_2_11 U2 (O[13], IN1[2], IN2);
  UB1BPPG_3_11 U3 (O[14], IN1[3], IN2);
  UB1BPPG_4_11 U4 (O[15], IN1[4], IN2);
  UB1BPPG_5_11 U5 (O[16], IN1[5], IN2);
  UB1BPPG_6_11 U6 (O[17], IN1[6], IN2);
  UB1BPPG_7_11 U7 (O[18], IN1[7], IN2);
  UB1BPPG_8_11 U8 (O[19], IN1[8], IN2);
  UB1BPPG_9_11 U9 (O[20], IN1[9], IN2);
  UB1BPPG_10_11 U10 (O[21], IN1[10], IN2);
  UB1BPPG_11_11 U11 (O[22], IN1[11], IN2);
  UB1BPPG_12_11 U12 (O[23], IN1[12], IN2);
  UB1BPPG_13_11 U13 (O[24], IN1[13], IN2);
  UB1BPPG_14_11 U14 (O[25], IN1[14], IN2);
  UB1BPPG_15_11 U15 (O[26], IN1[15], IN2);
endmodule

module UBVPPG_15_0_12 (O, IN1, IN2);
  output [27:12] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_12 U0 (O[12], IN1[0], IN2);
  UB1BPPG_1_12 U1 (O[13], IN1[1], IN2);
  UB1BPPG_2_12 U2 (O[14], IN1[2], IN2);
  UB1BPPG_3_12 U3 (O[15], IN1[3], IN2);
  UB1BPPG_4_12 U4 (O[16], IN1[4], IN2);
  UB1BPPG_5_12 U5 (O[17], IN1[5], IN2);
  UB1BPPG_6_12 U6 (O[18], IN1[6], IN2);
  UB1BPPG_7_12 U7 (O[19], IN1[7], IN2);
  UB1BPPG_8_12 U8 (O[20], IN1[8], IN2);
  UB1BPPG_9_12 U9 (O[21], IN1[9], IN2);
  UB1BPPG_10_12 U10 (O[22], IN1[10], IN2);
  UB1BPPG_11_12 U11 (O[23], IN1[11], IN2);
  UB1BPPG_12_12 U12 (O[24], IN1[12], IN2);
  UB1BPPG_13_12 U13 (O[25], IN1[13], IN2);
  UB1BPPG_14_12 U14 (O[26], IN1[14], IN2);
  UB1BPPG_15_12 U15 (O[27], IN1[15], IN2);
endmodule

module UBVPPG_15_0_13 (O, IN1, IN2);
  output [28:13] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_13 U0 (O[13], IN1[0], IN2);
  UB1BPPG_1_13 U1 (O[14], IN1[1], IN2);
  UB1BPPG_2_13 U2 (O[15], IN1[2], IN2);
  UB1BPPG_3_13 U3 (O[16], IN1[3], IN2);
  UB1BPPG_4_13 U4 (O[17], IN1[4], IN2);
  UB1BPPG_5_13 U5 (O[18], IN1[5], IN2);
  UB1BPPG_6_13 U6 (O[19], IN1[6], IN2);
  UB1BPPG_7_13 U7 (O[20], IN1[7], IN2);
  UB1BPPG_8_13 U8 (O[21], IN1[8], IN2);
  UB1BPPG_9_13 U9 (O[22], IN1[9], IN2);
  UB1BPPG_10_13 U10 (O[23], IN1[10], IN2);
  UB1BPPG_11_13 U11 (O[24], IN1[11], IN2);
  UB1BPPG_12_13 U12 (O[25], IN1[12], IN2);
  UB1BPPG_13_13 U13 (O[26], IN1[13], IN2);
  UB1BPPG_14_13 U14 (O[27], IN1[14], IN2);
  UB1BPPG_15_13 U15 (O[28], IN1[15], IN2);
endmodule

module UBVPPG_15_0_14 (O, IN1, IN2);
  output [29:14] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_14 U0 (O[14], IN1[0], IN2);
  UB1BPPG_1_14 U1 (O[15], IN1[1], IN2);
  UB1BPPG_2_14 U2 (O[16], IN1[2], IN2);
  UB1BPPG_3_14 U3 (O[17], IN1[3], IN2);
  UB1BPPG_4_14 U4 (O[18], IN1[4], IN2);
  UB1BPPG_5_14 U5 (O[19], IN1[5], IN2);
  UB1BPPG_6_14 U6 (O[20], IN1[6], IN2);
  UB1BPPG_7_14 U7 (O[21], IN1[7], IN2);
  UB1BPPG_8_14 U8 (O[22], IN1[8], IN2);
  UB1BPPG_9_14 U9 (O[23], IN1[9], IN2);
  UB1BPPG_10_14 U10 (O[24], IN1[10], IN2);
  UB1BPPG_11_14 U11 (O[25], IN1[11], IN2);
  UB1BPPG_12_14 U12 (O[26], IN1[12], IN2);
  UB1BPPG_13_14 U13 (O[27], IN1[13], IN2);
  UB1BPPG_14_14 U14 (O[28], IN1[14], IN2);
  UB1BPPG_15_14 U15 (O[29], IN1[15], IN2);
endmodule

module UBVPPG_15_0_15 (O, IN1, IN2);
  output [30:15] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_15 U0 (O[15], IN1[0], IN2);
  UB1BPPG_1_15 U1 (O[16], IN1[1], IN2);
  UB1BPPG_2_15 U2 (O[17], IN1[2], IN2);
  UB1BPPG_3_15 U3 (O[18], IN1[3], IN2);
  UB1BPPG_4_15 U4 (O[19], IN1[4], IN2);
  UB1BPPG_5_15 U5 (O[20], IN1[5], IN2);
  UB1BPPG_6_15 U6 (O[21], IN1[6], IN2);
  UB1BPPG_7_15 U7 (O[22], IN1[7], IN2);
  UB1BPPG_8_15 U8 (O[23], IN1[8], IN2);
  UB1BPPG_9_15 U9 (O[24], IN1[9], IN2);
  UB1BPPG_10_15 U10 (O[25], IN1[10], IN2);
  UB1BPPG_11_15 U11 (O[26], IN1[11], IN2);
  UB1BPPG_12_15 U12 (O[27], IN1[12], IN2);
  UB1BPPG_13_15 U13 (O[28], IN1[13], IN2);
  UB1BPPG_14_15 U14 (O[29], IN1[14], IN2);
  UB1BPPG_15_15 U15 (O[30], IN1[15], IN2);
endmodule

module UBVPPG_15_0_2 (O, IN1, IN2);
  output [17:2] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
  UB1BPPG_6_2 U6 (O[8], IN1[6], IN2);
  UB1BPPG_7_2 U7 (O[9], IN1[7], IN2);
  UB1BPPG_8_2 U8 (O[10], IN1[8], IN2);
  UB1BPPG_9_2 U9 (O[11], IN1[9], IN2);
  UB1BPPG_10_2 U10 (O[12], IN1[10], IN2);
  UB1BPPG_11_2 U11 (O[13], IN1[11], IN2);
  UB1BPPG_12_2 U12 (O[14], IN1[12], IN2);
  UB1BPPG_13_2 U13 (O[15], IN1[13], IN2);
  UB1BPPG_14_2 U14 (O[16], IN1[14], IN2);
  UB1BPPG_15_2 U15 (O[17], IN1[15], IN2);
endmodule

module UBVPPG_15_0_3 (O, IN1, IN2);
  output [18:3] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_3 U0 (O[3], IN1[0], IN2);
  UB1BPPG_1_3 U1 (O[4], IN1[1], IN2);
  UB1BPPG_2_3 U2 (O[5], IN1[2], IN2);
  UB1BPPG_3_3 U3 (O[6], IN1[3], IN2);
  UB1BPPG_4_3 U4 (O[7], IN1[4], IN2);
  UB1BPPG_5_3 U5 (O[8], IN1[5], IN2);
  UB1BPPG_6_3 U6 (O[9], IN1[6], IN2);
  UB1BPPG_7_3 U7 (O[10], IN1[7], IN2);
  UB1BPPG_8_3 U8 (O[11], IN1[8], IN2);
  UB1BPPG_9_3 U9 (O[12], IN1[9], IN2);
  UB1BPPG_10_3 U10 (O[13], IN1[10], IN2);
  UB1BPPG_11_3 U11 (O[14], IN1[11], IN2);
  UB1BPPG_12_3 U12 (O[15], IN1[12], IN2);
  UB1BPPG_13_3 U13 (O[16], IN1[13], IN2);
  UB1BPPG_14_3 U14 (O[17], IN1[14], IN2);
  UB1BPPG_15_3 U15 (O[18], IN1[15], IN2);
endmodule

module UBVPPG_15_0_4 (O, IN1, IN2);
  output [19:4] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
  UB1BPPG_6_4 U6 (O[10], IN1[6], IN2);
  UB1BPPG_7_4 U7 (O[11], IN1[7], IN2);
  UB1BPPG_8_4 U8 (O[12], IN1[8], IN2);
  UB1BPPG_9_4 U9 (O[13], IN1[9], IN2);
  UB1BPPG_10_4 U10 (O[14], IN1[10], IN2);
  UB1BPPG_11_4 U11 (O[15], IN1[11], IN2);
  UB1BPPG_12_4 U12 (O[16], IN1[12], IN2);
  UB1BPPG_13_4 U13 (O[17], IN1[13], IN2);
  UB1BPPG_14_4 U14 (O[18], IN1[14], IN2);
  UB1BPPG_15_4 U15 (O[19], IN1[15], IN2);
endmodule

module UBVPPG_15_0_5 (O, IN1, IN2);
  output [20:5] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_5 U0 (O[5], IN1[0], IN2);
  UB1BPPG_1_5 U1 (O[6], IN1[1], IN2);
  UB1BPPG_2_5 U2 (O[7], IN1[2], IN2);
  UB1BPPG_3_5 U3 (O[8], IN1[3], IN2);
  UB1BPPG_4_5 U4 (O[9], IN1[4], IN2);
  UB1BPPG_5_5 U5 (O[10], IN1[5], IN2);
  UB1BPPG_6_5 U6 (O[11], IN1[6], IN2);
  UB1BPPG_7_5 U7 (O[12], IN1[7], IN2);
  UB1BPPG_8_5 U8 (O[13], IN1[8], IN2);
  UB1BPPG_9_5 U9 (O[14], IN1[9], IN2);
  UB1BPPG_10_5 U10 (O[15], IN1[10], IN2);
  UB1BPPG_11_5 U11 (O[16], IN1[11], IN2);
  UB1BPPG_12_5 U12 (O[17], IN1[12], IN2);
  UB1BPPG_13_5 U13 (O[18], IN1[13], IN2);
  UB1BPPG_14_5 U14 (O[19], IN1[14], IN2);
  UB1BPPG_15_5 U15 (O[20], IN1[15], IN2);
endmodule

module UBVPPG_15_0_6 (O, IN1, IN2);
  output [21:6] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_6 U0 (O[6], IN1[0], IN2);
  UB1BPPG_1_6 U1 (O[7], IN1[1], IN2);
  UB1BPPG_2_6 U2 (O[8], IN1[2], IN2);
  UB1BPPG_3_6 U3 (O[9], IN1[3], IN2);
  UB1BPPG_4_6 U4 (O[10], IN1[4], IN2);
  UB1BPPG_5_6 U5 (O[11], IN1[5], IN2);
  UB1BPPG_6_6 U6 (O[12], IN1[6], IN2);
  UB1BPPG_7_6 U7 (O[13], IN1[7], IN2);
  UB1BPPG_8_6 U8 (O[14], IN1[8], IN2);
  UB1BPPG_9_6 U9 (O[15], IN1[9], IN2);
  UB1BPPG_10_6 U10 (O[16], IN1[10], IN2);
  UB1BPPG_11_6 U11 (O[17], IN1[11], IN2);
  UB1BPPG_12_6 U12 (O[18], IN1[12], IN2);
  UB1BPPG_13_6 U13 (O[19], IN1[13], IN2);
  UB1BPPG_14_6 U14 (O[20], IN1[14], IN2);
  UB1BPPG_15_6 U15 (O[21], IN1[15], IN2);
endmodule

module UBVPPG_15_0_7 (O, IN1, IN2);
  output [22:7] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_7 U0 (O[7], IN1[0], IN2);
  UB1BPPG_1_7 U1 (O[8], IN1[1], IN2);
  UB1BPPG_2_7 U2 (O[9], IN1[2], IN2);
  UB1BPPG_3_7 U3 (O[10], IN1[3], IN2);
  UB1BPPG_4_7 U4 (O[11], IN1[4], IN2);
  UB1BPPG_5_7 U5 (O[12], IN1[5], IN2);
  UB1BPPG_6_7 U6 (O[13], IN1[6], IN2);
  UB1BPPG_7_7 U7 (O[14], IN1[7], IN2);
  UB1BPPG_8_7 U8 (O[15], IN1[8], IN2);
  UB1BPPG_9_7 U9 (O[16], IN1[9], IN2);
  UB1BPPG_10_7 U10 (O[17], IN1[10], IN2);
  UB1BPPG_11_7 U11 (O[18], IN1[11], IN2);
  UB1BPPG_12_7 U12 (O[19], IN1[12], IN2);
  UB1BPPG_13_7 U13 (O[20], IN1[13], IN2);
  UB1BPPG_14_7 U14 (O[21], IN1[14], IN2);
  UB1BPPG_15_7 U15 (O[22], IN1[15], IN2);
endmodule

module UBVPPG_15_0_8 (O, IN1, IN2);
  output [23:8] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_8 U0 (O[8], IN1[0], IN2);
  UB1BPPG_1_8 U1 (O[9], IN1[1], IN2);
  UB1BPPG_2_8 U2 (O[10], IN1[2], IN2);
  UB1BPPG_3_8 U3 (O[11], IN1[3], IN2);
  UB1BPPG_4_8 U4 (O[12], IN1[4], IN2);
  UB1BPPG_5_8 U5 (O[13], IN1[5], IN2);
  UB1BPPG_6_8 U6 (O[14], IN1[6], IN2);
  UB1BPPG_7_8 U7 (O[15], IN1[7], IN2);
  UB1BPPG_8_8 U8 (O[16], IN1[8], IN2);
  UB1BPPG_9_8 U9 (O[17], IN1[9], IN2);
  UB1BPPG_10_8 U10 (O[18], IN1[10], IN2);
  UB1BPPG_11_8 U11 (O[19], IN1[11], IN2);
  UB1BPPG_12_8 U12 (O[20], IN1[12], IN2);
  UB1BPPG_13_8 U13 (O[21], IN1[13], IN2);
  UB1BPPG_14_8 U14 (O[22], IN1[14], IN2);
  UB1BPPG_15_8 U15 (O[23], IN1[15], IN2);
endmodule

module UBVPPG_15_0_9 (O, IN1, IN2);
  output [24:9] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_9 U0 (O[9], IN1[0], IN2);
  UB1BPPG_1_9 U1 (O[10], IN1[1], IN2);
  UB1BPPG_2_9 U2 (O[11], IN1[2], IN2);
  UB1BPPG_3_9 U3 (O[12], IN1[3], IN2);
  UB1BPPG_4_9 U4 (O[13], IN1[4], IN2);
  UB1BPPG_5_9 U5 (O[14], IN1[5], IN2);
  UB1BPPG_6_9 U6 (O[15], IN1[6], IN2);
  UB1BPPG_7_9 U7 (O[16], IN1[7], IN2);
  UB1BPPG_8_9 U8 (O[17], IN1[8], IN2);
  UB1BPPG_9_9 U9 (O[18], IN1[9], IN2);
  UB1BPPG_10_9 U10 (O[19], IN1[10], IN2);
  UB1BPPG_11_9 U11 (O[20], IN1[11], IN2);
  UB1BPPG_12_9 U12 (O[21], IN1[12], IN2);
  UB1BPPG_13_9 U13 (O[22], IN1[13], IN2);
  UB1BPPG_14_9 U14 (O[23], IN1[14], IN2);
  UB1BPPG_15_9 U15 (O[24], IN1[15], IN2);
endmodule

