/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: Multiplier_14_0_1000

  Number system: Unsigned binary
  Multiplicand length: 15
  Multiplier length: 15
  Partial product generation: Simple PPG
  Partial product accumulation: Redundant binary addition tree
  Final stage addition: Carry-skip adder (fixed-block-size)
----------------------------------------------------------------------------*/

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module SignP_0(O);
  output O;
  assign O = 0;
endmodule

module BWCPN_1(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_2(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_3(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_4(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_5(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_6(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_7(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_8(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_9(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_10(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_11(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_12(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_13(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_14(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_15(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module NUBBBG_1(O, S);
  output O;
  input S;
  assign O = ~ S;
endmodule

module UBHBBG_16(O, S);
  output O;
  input S;
  assign O = ~ S;
endmodule

module UB1DCON_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_15_15(O);
  output [15:15] O;
  assign O[15] = 0;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUBZero_16_16(O);
  output [16:16] O;
  assign O[16] = 0;
endmodule

module NUBZero_0_0(O);
  output [0:0] O;
  assign O[0] = 0;
endmodule

module NUB1DCON_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module SD2DigitCom_0(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_1(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_2(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_3(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_4(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_5(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_6(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_7(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_8(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_9(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_10(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_11(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_12(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_13(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_14(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_15(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_16(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module BWCPN_16(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_17(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module NUBBBG_3(O, S);
  output O;
  input S;
  assign O = ~ S;
endmodule

module UBHBBG_18(O, S);
  output O;
  input S;
  assign O = ~ S;
endmodule

module UB1DCON_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_17_17(O);
  output [17:17] O;
  assign O[17] = 0;
endmodule

module UB1DCON_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUBZero_18_18(O);
  output [18:18] O;
  assign O[18] = 0;
endmodule

module NUBZero_2_2(O);
  output [2:2] O;
  assign O[2] = 0;
endmodule

module NUB1DCON_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module SD2DigitCom_17(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_18(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module BWCPN_18(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_19(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module NUBBBG_5(O, S);
  output O;
  input S;
  assign O = ~ S;
endmodule

module UBHBBG_20(O, S);
  output O;
  input S;
  assign O = ~ S;
endmodule

module UB1DCON_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_19_19(O);
  output [19:19] O;
  assign O[19] = 0;
endmodule

module UB1DCON_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUBZero_20_20(O);
  output [20:20] O;
  assign O[20] = 0;
endmodule

module NUBZero_4_4(O);
  output [4:4] O;
  assign O[4] = 0;
endmodule

module NUB1DCON_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module SD2DigitCom_19(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_20(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module UB1BPPG_0_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module BWCPN_20(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_21(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module NUBBBG_7(O, S);
  output O;
  input S;
  assign O = ~ S;
endmodule

module UBHBBG_22(O, S);
  output O;
  input S;
  assign O = ~ S;
endmodule

module UB1DCON_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_21_21(O);
  output [21:21] O;
  assign O[21] = 0;
endmodule

module UB1DCON_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUBZero_22_22(O);
  output [22:22] O;
  assign O[22] = 0;
endmodule

module NUBZero_6_6(O);
  output [6:6] O;
  assign O[6] = 0;
endmodule

module NUB1DCON_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_21(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module SD2DigitCom_21(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_22(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module UB1BPPG_0_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module BWCPN_22(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_23(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module NUBBBG_9(O, S);
  output O;
  input S;
  assign O = ~ S;
endmodule

module UBHBBG_24(O, S);
  output O;
  input S;
  assign O = ~ S;
endmodule

module UB1DCON_24(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_23_23(O);
  output [23:23] O;
  assign O[23] = 0;
endmodule

module UB1DCON_21(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUBZero_24_24(O);
  output [24:24] O;
  assign O[24] = 0;
endmodule

module NUBZero_8_8(O);
  output [8:8] O;
  assign O[8] = 0;
endmodule

module NUB1DCON_24(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_23(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module SD2DigitCom_23(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_24(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module UB1BPPG_0_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module BWCPN_24(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_25(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module NUBBBG_11(O, S);
  output O;
  input S;
  assign O = ~ S;
endmodule

module UBHBBG_26(O, S);
  output O;
  input S;
  assign O = ~ S;
endmodule

module UB1DCON_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_25_25(O);
  output [25:25] O;
  assign O[25] = 0;
endmodule

module UB1DCON_23(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUBZero_26_26(O);
  output [26:26] O;
  assign O[26] = 0;
endmodule

module NUBZero_10_10(O);
  output [10:10] O;
  assign O[10] = 0;
endmodule

module NUB1DCON_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_25(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module SD2DigitCom_25(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_26(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module UB1BPPG_0_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module BWCPN_26(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module BWCPN_27(O, I, S);
  output O;
  input I;
  input S;
  assign O = S ^ ( ~ I );
endmodule

module NUBBBG_13(O, S);
  output O;
  input S;
  assign O = ~ S;
endmodule

module UBHBBG_28(O, S);
  output O;
  input S;
  assign O = ~ S;
endmodule

module UB1DCON_28(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_27_27(O);
  output [27:27] O;
  assign O[27] = 0;
endmodule

module UB1DCON_25(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUBZero_28_28(O);
  output [28:28] O;
  assign O[28] = 0;
endmodule

module NUBZero_12_12(O);
  output [12:12] O;
  assign O[12] = 0;
endmodule

module NUB1DCON_28(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module NUB1DCON_27(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module SD2DigitCom_27(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitCom_28(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module UB1BPPG_0_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBZero_28_14(O);
  output [28:14] O;
  assign O[14] = 0;
  assign O[15] = 0;
  assign O[16] = 0;
  assign O[17] = 0;
  assign O[18] = 0;
  assign O[19] = 0;
  assign O[20] = 0;
  assign O[21] = 0;
  assign O[22] = 0;
  assign O[23] = 0;
  assign O[24] = 0;
  assign O[25] = 0;
  assign O[26] = 0;
  assign O[27] = 0;
  assign O[28] = 0;
endmodule

module UBZero_13_1(O);
  output [13:1] O;
  assign O[1] = 0;
  assign O[2] = 0;
  assign O[3] = 0;
  assign O[4] = 0;
  assign O[5] = 0;
  assign O[6] = 0;
  assign O[7] = 0;
  assign O[8] = 0;
  assign O[9] = 0;
  assign O[10] = 0;
  assign O[11] = 0;
  assign O[12] = 0;
  assign O[13] = 0;
endmodule

module UB1DCON_27(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module SD2_PN_A_Zero_18_000(O_p, O_n);
  output [18:17] O_p, O_n;
  assign O_p[17] = 0;
  assign O_n[17] = 0;
  assign O_p[18] = 0;
  assign O_n[18] = 0;
endmodule

module SD2_PN_A1DCON_17(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_18(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_0(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_1(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_2(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_3(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_4(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_5(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_6(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_7(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_8(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_9(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_10(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_11(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_12(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_13(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_14(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_15(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_16(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module UBZero_2_2(O);
  output [2:2] O;
  assign O[2] = 0;
endmodule

module SD2DigitDecom_PN_000(X, Y, I_p, I_n);
  output [2:2] X;
  output [2:2] Y;
  input [2:2] I_p, I_n;
  assign X = ~ I_n[2];
  assign Y = I_p[2];
endmodule

module UBFA_2(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_3(O, I);
  output [3:3] O;
  input [3:3] I;
  assign O[3] = ~ I[3];
endmodule

module SD2DigitDecom_PN_001(X, Y, I_p, I_n);
  output [3:3] X;
  output [3:3] Y;
  input [3:3] I_p, I_n;
  assign X = ~ I_n[3];
  assign Y = I_p[3];
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_4(O, I);
  output [4:4] O;
  input [4:4] I;
  assign O[4] = ~ I[4];
endmodule

module SD2DigitDecom_PN_002(X, Y, I_p, I_n);
  output [4:4] X;
  output [4:4] Y;
  input [4:4] I_p, I_n;
  assign X = ~ I_n[4];
  assign Y = I_p[4];
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_5(O, I);
  output [5:5] O;
  input [5:5] I;
  assign O[5] = ~ I[5];
endmodule

module SD2DigitDecom_PN_003(X, Y, I_p, I_n);
  output [5:5] X;
  output [5:5] Y;
  input [5:5] I_p, I_n;
  assign X = ~ I_n[5];
  assign Y = I_p[5];
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_6(O, I);
  output [6:6] O;
  input [6:6] I;
  assign O[6] = ~ I[6];
endmodule

module SD2DigitDecom_PN_004(X, Y, I_p, I_n);
  output [6:6] X;
  output [6:6] Y;
  input [6:6] I_p, I_n;
  assign X = ~ I_n[6];
  assign Y = I_p[6];
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_7(O, I);
  output [7:7] O;
  input [7:7] I;
  assign O[7] = ~ I[7];
endmodule

module SD2DigitDecom_PN_005(X, Y, I_p, I_n);
  output [7:7] X;
  output [7:7] Y;
  input [7:7] I_p, I_n;
  assign X = ~ I_n[7];
  assign Y = I_p[7];
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_8(O, I);
  output [8:8] O;
  input [8:8] I;
  assign O[8] = ~ I[8];
endmodule

module SD2DigitDecom_PN_006(X, Y, I_p, I_n);
  output [8:8] X;
  output [8:8] Y;
  input [8:8] I_p, I_n;
  assign X = ~ I_n[8];
  assign Y = I_p[8];
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_9(O, I);
  output [9:9] O;
  input [9:9] I;
  assign O[9] = ~ I[9];
endmodule

module SD2DigitDecom_PN_007(X, Y, I_p, I_n);
  output [9:9] X;
  output [9:9] Y;
  input [9:9] I_p, I_n;
  assign X = ~ I_n[9];
  assign Y = I_p[9];
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_10(O, I);
  output [10:10] O;
  input [10:10] I;
  assign O[10] = ~ I[10];
endmodule

module SD2DigitDecom_PN_008(X, Y, I_p, I_n);
  output [10:10] X;
  output [10:10] Y;
  input [10:10] I_p, I_n;
  assign X = ~ I_n[10];
  assign Y = I_p[10];
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_11(O, I);
  output [11:11] O;
  input [11:11] I;
  assign O[11] = ~ I[11];
endmodule

module SD2DigitDecom_PN_009(X, Y, I_p, I_n);
  output [11:11] X;
  output [11:11] Y;
  input [11:11] I_p, I_n;
  assign X = ~ I_n[11];
  assign Y = I_p[11];
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_12(O, I);
  output [12:12] O;
  input [12:12] I;
  assign O[12] = ~ I[12];
endmodule

module SD2DigitDecom_PN_010(X, Y, I_p, I_n);
  output [12:12] X;
  output [12:12] Y;
  input [12:12] I_p, I_n;
  assign X = ~ I_n[12];
  assign Y = I_p[12];
endmodule

module UBFA_12(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_13(O, I);
  output [13:13] O;
  input [13:13] I;
  assign O[13] = ~ I[13];
endmodule

module SD2DigitDecom_PN_011(X, Y, I_p, I_n);
  output [13:13] X;
  output [13:13] Y;
  input [13:13] I_p, I_n;
  assign X = ~ I_n[13];
  assign Y = I_p[13];
endmodule

module UBFA_13(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_14(O, I);
  output [14:14] O;
  input [14:14] I;
  assign O[14] = ~ I[14];
endmodule

module SD2DigitDecom_PN_012(X, Y, I_p, I_n);
  output [14:14] X;
  output [14:14] Y;
  input [14:14] I_p, I_n;
  assign X = ~ I_n[14];
  assign Y = I_p[14];
endmodule

module UBFA_14(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_15(O, I);
  output [15:15] O;
  input [15:15] I;
  assign O[15] = ~ I[15];
endmodule

module SD2DigitDecom_PN_013(X, Y, I_p, I_n);
  output [15:15] X;
  output [15:15] Y;
  input [15:15] I_p, I_n;
  assign X = ~ I_n[15];
  assign Y = I_p[15];
endmodule

module UBFA_15(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_16(O, I);
  output [16:16] O;
  input [16:16] I;
  assign O[16] = ~ I[16];
endmodule

module SD2DigitDecom_PN_014(X, Y, I_p, I_n);
  output [16:16] X;
  output [16:16] Y;
  input [16:16] I_p, I_n;
  assign X = ~ I_n[16];
  assign Y = I_p[16];
endmodule

module UBFA_16(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_17(O, I);
  output [17:17] O;
  input [17:17] I;
  assign O[17] = ~ I[17];
endmodule

module SD2DigitDecom_PN_015(X, Y, I_p, I_n);
  output [17:17] X;
  output [17:17] Y;
  input [17:17] I_p, I_n;
  assign X = ~ I_n[17];
  assign Y = I_p[17];
endmodule

module UBFA_17(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_18(O, I);
  output [18:18] O;
  input [18:18] I;
  assign O[18] = ~ I[18];
endmodule

module SD2DigitDecom_PN_016(X, Y, I_p, I_n);
  output [18:18] X;
  output [18:18] Y;
  input [18:18] I_p, I_n;
  assign X = ~ I_n[18];
  assign Y = I_p[18];
endmodule

module UBFA_18(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_19(O, I);
  output [19:19] O;
  input [19:19] I;
  assign O[19] = ~ I[19];
endmodule

module SD2_PN_A_Zero_22_000(O_p, O_n);
  output [22:21] O_p, O_n;
  assign O_p[21] = 0;
  assign O_n[21] = 0;
  assign O_p[22] = 0;
  assign O_n[22] = 0;
endmodule

module SD2_PN_A1DCON_21(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_22(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_19(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_20(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module UBZero_6_6(O);
  output [6:6] O;
  assign O[6] = 0;
endmodule

module SD2DigitDecom_PN_017(X, Y, I_p, I_n);
  output [19:19] X;
  output [19:19] Y;
  input [19:19] I_p, I_n;
  assign X = ~ I_n[19];
  assign Y = I_p[19];
endmodule

module UBFA_19(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_20(O, I);
  output [20:20] O;
  input [20:20] I;
  assign O[20] = ~ I[20];
endmodule

module SD2DigitDecom_PN_018(X, Y, I_p, I_n);
  output [20:20] X;
  output [20:20] Y;
  input [20:20] I_p, I_n;
  assign X = ~ I_n[20];
  assign Y = I_p[20];
endmodule

module UBFA_20(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_21(O, I);
  output [21:21] O;
  input [21:21] I;
  assign O[21] = ~ I[21];
endmodule

module SD2DigitDecom_PN_019(X, Y, I_p, I_n);
  output [21:21] X;
  output [21:21] Y;
  input [21:21] I_p, I_n;
  assign X = ~ I_n[21];
  assign Y = I_p[21];
endmodule

module UBFA_21(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_22(O, I);
  output [22:22] O;
  input [22:22] I;
  assign O[22] = ~ I[22];
endmodule

module SD2DigitDecom_PN_020(X, Y, I_p, I_n);
  output [22:22] X;
  output [22:22] Y;
  input [22:22] I_p, I_n;
  assign X = ~ I_n[22];
  assign Y = I_p[22];
endmodule

module UBFA_22(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_23(O, I);
  output [23:23] O;
  input [23:23] I;
  assign O[23] = ~ I[23];
endmodule

module SD2_PN_A_Zero_26_000(O_p, O_n);
  output [26:25] O_p, O_n;
  assign O_p[25] = 0;
  assign O_n[25] = 0;
  assign O_p[26] = 0;
  assign O_n[26] = 0;
endmodule

module SD2_PN_A1DCON_25(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_26(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_23(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_24(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module UBZero_10_10(O);
  output [10:10] O;
  assign O[10] = 0;
endmodule

module SD2DigitDecom_PN_021(X, Y, I_p, I_n);
  output [23:23] X;
  output [23:23] Y;
  input [23:23] I_p, I_n;
  assign X = ~ I_n[23];
  assign Y = I_p[23];
endmodule

module UBFA_23(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_24(O, I);
  output [24:24] O;
  input [24:24] I;
  assign O[24] = ~ I[24];
endmodule

module SD2DigitDecom_PN_022(X, Y, I_p, I_n);
  output [24:24] X;
  output [24:24] Y;
  input [24:24] I_p, I_n;
  assign X = ~ I_n[24];
  assign Y = I_p[24];
endmodule

module UBFA_24(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_25(O, I);
  output [25:25] O;
  input [25:25] I;
  assign O[25] = ~ I[25];
endmodule

module SD2DigitDecom_PN_023(X, Y, I_p, I_n);
  output [25:25] X;
  output [25:25] Y;
  input [25:25] I_p, I_n;
  assign X = ~ I_n[25];
  assign Y = I_p[25];
endmodule

module UBFA_25(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_26(O, I);
  output [26:26] O;
  input [26:26] I;
  assign O[26] = ~ I[26];
endmodule

module SD2DigitDecom_PN_024(X, Y, I_p, I_n);
  output [26:26] X;
  output [26:26] Y;
  input [26:26] I_p, I_n;
  assign X = ~ I_n[26];
  assign Y = I_p[26];
endmodule

module UBFA_26(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_27(O, I);
  output [27:27] O;
  input [27:27] I;
  assign O[27] = ~ I[27];
endmodule

module UBZero_12_12(O);
  output [12:12] O;
  assign O[12] = 0;
endmodule

module SD2DigitDecom_PN_025(X, Y, I_p, I_n);
  output [27:27] X;
  output [27:27] Y;
  input [27:27] I_p, I_n;
  assign X = ~ I_n[27];
  assign Y = I_p[27];
endmodule

module UBFA_27(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_28(O, I);
  output [28:28] O;
  input [28:28] I;
  assign O[28] = ~ I[28];
endmodule

module SD2DigitDecom_PN_026(X, Y, I_p, I_n);
  output [28:28] X;
  output [28:28] Y;
  input [28:28] I_p, I_n;
  assign X = ~ I_n[28];
  assign Y = I_p[28];
endmodule

module UBFA_28(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_29(O, I);
  output [29:29] O;
  input [29:29] I;
  assign O[29] = ~ I[29];
endmodule

module SD2DigitCom_29(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A_Zero_23_000(O_p, O_n);
  output [23:20] O_p, O_n;
  assign O_p[20] = 0;
  assign O_n[20] = 0;
  assign O_p[21] = 0;
  assign O_n[21] = 0;
  assign O_p[22] = 0;
  assign O_n[22] = 0;
  assign O_p[23] = 0;
  assign O_n[23] = 0;
endmodule

module UBZero_4_4(O);
  output [4:4] O;
  assign O[4] = 0;
endmodule

module SD2_PN_A_Zero_29_000(O_p, O_n);
  output [29:28] O_p, O_n;
  assign O_p[28] = 0;
  assign O_n[28] = 0;
  assign O_p[29] = 0;
  assign O_n[29] = 0;
endmodule

module SD2_PN_A1DCON_28(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_29(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A1DCON_27(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module UBZero_8_8(O);
  output [8:8] O;
  assign O[8] = 0;
endmodule

module SD2DigitDecom_PN_027(X, Y, I_p, I_n);
  output [29:29] X;
  output [29:29] Y;
  input [29:29] I_p, I_n;
  assign X = ~ I_n[29];
  assign Y = I_p[29];
endmodule

module UBFA_29(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_30(O, I);
  output [30:30] O;
  input [30:30] I;
  assign O[30] = ~ I[30];
endmodule

module SD2DigitCom_30(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2_PN_A_Zero_30_000(O_p, O_n);
  output [30:25] O_p, O_n;
  assign O_p[25] = 0;
  assign O_n[25] = 0;
  assign O_p[26] = 0;
  assign O_n[26] = 0;
  assign O_p[27] = 0;
  assign O_n[27] = 0;
  assign O_p[28] = 0;
  assign O_n[28] = 0;
  assign O_p[29] = 0;
  assign O_n[29] = 0;
  assign O_p[30] = 0;
  assign O_n[30] = 0;
endmodule

module SD2_PN_A1DCON_30(O_p, O_n, I_p, I_n);
  output O_p, O_n;
  input I_p, I_n;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module UBZero_1_1(O);
  output [1:1] O;
  assign O[1] = 0;
endmodule

module NUBZero_1_1(O);
  output [1:1] O;
  assign O[1] = 0;
endmodule

module SD2DigitDecom_PN_028(X, Y, I_p, I_n);
  output [1:1] X;
  output [1:1] Y;
  input [1:1] I_p, I_n;
  assign X = ~ I_n[1];
  assign Y = I_p[1];
endmodule

module UBFA_1(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_2(O, I);
  output [2:2] O;
  input [2:2] I;
  assign O[2] = ~ I[2];
endmodule

module SD2DigitDecom_PN_029(X, Y, I_p, I_n);
  output [30:30] X;
  output [30:30] Y;
  input [30:30] I_p, I_n;
  assign X = ~ I_n[30];
  assign Y = I_p[30];
endmodule

module UBFA_30(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBInv_31(O, I);
  output [31:31] O;
  input [31:31] I;
  assign O[31] = ~ I[31];
endmodule

module SD2DigitCom_31(O_p, O_n, I_n, I_p);
  output O_p, O_n;
  input I_n;
  input I_p;
  assign O_p = I_p;
  assign O_n = I_n;
endmodule

module SD2DigitDecom_PN_030(X, Y, I_p, I_n);
  output [0:0] X;
  output [0:0] Y;
  input [0:0] I_p, I_n;
  assign X = ~ I_n[0];
  assign Y = I_p[0];
endmodule

module SD2DigitDecom_PN_031(X, Y, I_p, I_n);
  output [31:31] X;
  output [31:31] Y;
  input [31:31] I_p, I_n;
  assign X = ~ I_n[31];
  assign Y = I_p[31];
endmodule

module UBOne_0(O);
  output O;
  assign O = 1;
endmodule

module UBHA_0(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_0(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_0 U0 (C_0, S_0, X, Y);
  UBHA_0 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_1(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_1(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_1 U0 (C_0, S_0, X, Y);
  UBHA_1 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_2(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_2 U0 (C_0, S_0, X, Y);
  UBHA_2 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_3(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_3 U0 (C_0, S_0, X, Y);
  UBHA_3 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_3_0(Co, S, X, Y, Ci);
  output Co;
  output [3:0] S;
  input Ci;
  input [3:0] X;
  input [3:0] Y;
  wire C1;
  wire C2;
  wire C3;
  wire C4;
  wire P0;
  wire P1;
  wire P2;
  wire P3;
  wire Sk;
  assign Sk = ( P0 & P1 & P2 & P3 ) & Ci;
  assign Co = C4 | Sk;
  UBPFA_0 U0 (C1, S[0], P0, X[0], Y[0], Ci);
  UBPFA_1 U1 (C2, S[1], P1, X[1], Y[1], C1);
  UBPFA_2 U2 (C3, S[2], P2, X[2], Y[2], C2);
  UBPFA_3 U3 (C4, S[3], P3, X[3], Y[3], C3);
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_4(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_4 U0 (C_0, S_0, X, Y);
  UBHA_4 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_5(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_5(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_5 U0 (C_0, S_0, X, Y);
  UBHA_5 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_6(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_6(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_6 U0 (C_0, S_0, X, Y);
  UBHA_6 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_7(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_7(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_7 U0 (C_0, S_0, X, Y);
  UBHA_7 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_7_4(Co, S, X, Y, Ci);
  output Co;
  output [7:4] S;
  input Ci;
  input [7:4] X;
  input [7:4] Y;
  wire C5;
  wire C6;
  wire C7;
  wire C8;
  wire P4;
  wire P5;
  wire P6;
  wire P7;
  wire Sk;
  assign Sk = ( P4 & P5 & P6 & P7 ) & Ci;
  assign Co = C8 | Sk;
  UBPFA_4 U0 (C5, S[4], P4, X[4], Y[4], Ci);
  UBPFA_5 U1 (C6, S[5], P5, X[5], Y[5], C5);
  UBPFA_6 U2 (C7, S[6], P6, X[6], Y[6], C6);
  UBPFA_7 U3 (C8, S[7], P7, X[7], Y[7], C7);
endmodule

module UBHA_8(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_8(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_8 U0 (C_0, S_0, X, Y);
  UBHA_8 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_9(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_9(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_9 U0 (C_0, S_0, X, Y);
  UBHA_9 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_10(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_10(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_10 U0 (C_0, S_0, X, Y);
  UBHA_10 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_11(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_11(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_11 U0 (C_0, S_0, X, Y);
  UBHA_11 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_11_8(Co, S, X, Y, Ci);
  output Co;
  output [11:8] S;
  input Ci;
  input [11:8] X;
  input [11:8] Y;
  wire C10;
  wire C11;
  wire C12;
  wire C9;
  wire P10;
  wire P11;
  wire P8;
  wire P9;
  wire Sk;
  assign Sk = ( P8 & P9 & P10 & P11 ) & Ci;
  assign Co = C12 | Sk;
  UBPFA_8 U0 (C9, S[8], P8, X[8], Y[8], Ci);
  UBPFA_9 U1 (C10, S[9], P9, X[9], Y[9], C9);
  UBPFA_10 U2 (C11, S[10], P10, X[10], Y[10], C10);
  UBPFA_11 U3 (C12, S[11], P11, X[11], Y[11], C11);
endmodule

module UBHA_12(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_12(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_12 U0 (C_0, S_0, X, Y);
  UBHA_12 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_13(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_13(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_13 U0 (C_0, S_0, X, Y);
  UBHA_13 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_14(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_14(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_14 U0 (C_0, S_0, X, Y);
  UBHA_14 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_15(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_15(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_15 U0 (C_0, S_0, X, Y);
  UBHA_15 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_15_12(Co, S, X, Y, Ci);
  output Co;
  output [15:12] S;
  input Ci;
  input [15:12] X;
  input [15:12] Y;
  wire C13;
  wire C14;
  wire C15;
  wire C16;
  wire P12;
  wire P13;
  wire P14;
  wire P15;
  wire Sk;
  assign Sk = ( P12 & P13 & P14 & P15 ) & Ci;
  assign Co = C16 | Sk;
  UBPFA_12 U0 (C13, S[12], P12, X[12], Y[12], Ci);
  UBPFA_13 U1 (C14, S[13], P13, X[13], Y[13], C13);
  UBPFA_14 U2 (C15, S[14], P14, X[14], Y[14], C14);
  UBPFA_15 U3 (C16, S[15], P15, X[15], Y[15], C15);
endmodule

module UBHA_16(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_16(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_16 U0 (C_0, S_0, X, Y);
  UBHA_16 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_17(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_17(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_17 U0 (C_0, S_0, X, Y);
  UBHA_17 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_18(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_18(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_18 U0 (C_0, S_0, X, Y);
  UBHA_18 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_19(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_19(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_19 U0 (C_0, S_0, X, Y);
  UBHA_19 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_19_16(Co, S, X, Y, Ci);
  output Co;
  output [19:16] S;
  input Ci;
  input [19:16] X;
  input [19:16] Y;
  wire C17;
  wire C18;
  wire C19;
  wire C20;
  wire P16;
  wire P17;
  wire P18;
  wire P19;
  wire Sk;
  assign Sk = ( P16 & P17 & P18 & P19 ) & Ci;
  assign Co = C20 | Sk;
  UBPFA_16 U0 (C17, S[16], P16, X[16], Y[16], Ci);
  UBPFA_17 U1 (C18, S[17], P17, X[17], Y[17], C17);
  UBPFA_18 U2 (C19, S[18], P18, X[18], Y[18], C18);
  UBPFA_19 U3 (C20, S[19], P19, X[19], Y[19], C19);
endmodule

module UBHA_20(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_20(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_20 U0 (C_0, S_0, X, Y);
  UBHA_20 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_21(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_21(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_21 U0 (C_0, S_0, X, Y);
  UBHA_21 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_22(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_22(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_22 U0 (C_0, S_0, X, Y);
  UBHA_22 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_23(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_23(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_23 U0 (C_0, S_0, X, Y);
  UBHA_23 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_23_20(Co, S, X, Y, Ci);
  output Co;
  output [23:20] S;
  input Ci;
  input [23:20] X;
  input [23:20] Y;
  wire C21;
  wire C22;
  wire C23;
  wire C24;
  wire P20;
  wire P21;
  wire P22;
  wire P23;
  wire Sk;
  assign Sk = ( P20 & P21 & P22 & P23 ) & Ci;
  assign Co = C24 | Sk;
  UBPFA_20 U0 (C21, S[20], P20, X[20], Y[20], Ci);
  UBPFA_21 U1 (C22, S[21], P21, X[21], Y[21], C21);
  UBPFA_22 U2 (C23, S[22], P22, X[22], Y[22], C22);
  UBPFA_23 U3 (C24, S[23], P23, X[23], Y[23], C23);
endmodule

module UBHA_24(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_24(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_24 U0 (C_0, S_0, X, Y);
  UBHA_24 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_25(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_25(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_25 U0 (C_0, S_0, X, Y);
  UBHA_25 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_26(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_26(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_26 U0 (C_0, S_0, X, Y);
  UBHA_26 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_27(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_27(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_27 U0 (C_0, S_0, X, Y);
  UBHA_27 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_27_24(Co, S, X, Y, Ci);
  output Co;
  output [27:24] S;
  input Ci;
  input [27:24] X;
  input [27:24] Y;
  wire C25;
  wire C26;
  wire C27;
  wire C28;
  wire P24;
  wire P25;
  wire P26;
  wire P27;
  wire Sk;
  assign Sk = ( P24 & P25 & P26 & P27 ) & Ci;
  assign Co = C28 | Sk;
  UBPFA_24 U0 (C25, S[24], P24, X[24], Y[24], Ci);
  UBPFA_25 U1 (C26, S[25], P25, X[25], Y[25], C25);
  UBPFA_26 U2 (C27, S[26], P26, X[26], Y[26], C26);
  UBPFA_27 U3 (C28, S[27], P27, X[27], Y[27], C27);
endmodule

module UBHA_28(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_28(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_28 U0 (C_0, S_0, X, Y);
  UBHA_28 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_29(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_29(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_29 U0 (C_0, S_0, X, Y);
  UBHA_29 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_30(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_30(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_30 U0 (C_0, S_0, X, Y);
  UBHA_30 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_31(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_31(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_31 U0 (C_0, S_0, X, Y);
  UBHA_31 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_31_28(Co, S, X, Y, Ci);
  output Co;
  output [31:28] S;
  input Ci;
  input [31:28] X;
  input [31:28] Y;
  wire C29;
  wire C30;
  wire C31;
  wire C32;
  wire P28;
  wire P29;
  wire P30;
  wire P31;
  wire Sk;
  assign Sk = ( P28 & P29 & P30 & P31 ) & Ci;
  assign Co = C32 | Sk;
  UBPFA_28 U0 (C29, S[28], P28, X[28], Y[28], Ci);
  UBPFA_29 U1 (C30, S[29], P29, X[29], Y[29], C29);
  UBPFA_30 U2 (C31, S[30], P30, X[30], Y[30], C30);
  UBPFA_31 U3 (C32, S[31], P31, X[31], Y[31], C31);
endmodule

module UBPriFCSkA_31_0(S, X, Y, Cin);
  output [32:0] S;
  input Cin;
  input [31:0] X;
  input [31:0] Y;
  wire C12;
  wire C16;
  wire C20;
  wire C24;
  wire C28;
  wire C4;
  wire C8;
  UBCSkB_3_0 U0 (C4, S[3:0], X[3:0], Y[3:0], Cin);
  UBCSkB_7_4 U1 (C8, S[7:4], X[7:4], Y[7:4], C4);
  UBCSkB_11_8 U2 (C12, S[11:8], X[11:8], Y[11:8], C8);
  UBCSkB_15_12 U3 (C16, S[15:12], X[15:12], Y[15:12], C12);
  UBCSkB_19_16 U4 (C20, S[19:16], X[19:16], Y[19:16], C16);
  UBCSkB_23_20 U5 (C24, S[23:20], X[23:20], Y[23:20], C20);
  UBCSkB_27_24 U6 (C28, S[27:24], X[27:24], Y[27:24], C24);
  UBCSkB_31_28 U7 (S[32], S[31:28], X[31:28], Y[31:28], C28);
endmodule

module UBInv_32(O, I);
  output [32:32] O;
  input [32:32] I;
  assign O[32] = ~ I[32];
endmodule

module TCCom_32_0(O, I1, I2);
  output [32:0] O;
  input [32:32] I1;
  input [31:0] I2;
  assign O[32] = I1;
  assign O[0] = I2[0];
  assign O[1] = I2[1];
  assign O[2] = I2[2];
  assign O[3] = I2[3];
  assign O[4] = I2[4];
  assign O[5] = I2[5];
  assign O[6] = I2[6];
  assign O[7] = I2[7];
  assign O[8] = I2[8];
  assign O[9] = I2[9];
  assign O[10] = I2[10];
  assign O[11] = I2[11];
  assign O[12] = I2[12];
  assign O[13] = I2[13];
  assign O[14] = I2[14];
  assign O[15] = I2[15];
  assign O[16] = I2[16];
  assign O[17] = I2[17];
  assign O[18] = I2[18];
  assign O[19] = I2[19];
  assign O[20] = I2[20];
  assign O[21] = I2[21];
  assign O[22] = I2[22];
  assign O[23] = I2[23];
  assign O[24] = I2[24];
  assign O[25] = I2[25];
  assign O[26] = I2[26];
  assign O[27] = I2[27];
  assign O[28] = I2[28];
  assign O[29] = I2[29];
  assign O[30] = I2[30];
  assign O[31] = I2[31];
endmodule

module Multiplier_14_0_1000(P, IN1, IN2);
  output [29:0] P;
  input [14:0] IN1;
  input [14:0] IN2;
  wire [32:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  assign P[12] = W[12];
  assign P[13] = W[13];
  assign P[14] = W[14];
  assign P[15] = W[15];
  assign P[16] = W[16];
  assign P[17] = W[17];
  assign P[18] = W[18];
  assign P[19] = W[19];
  assign P[20] = W[20];
  assign P[21] = W[21];
  assign P[22] = W[22];
  assign P[23] = W[23];
  assign P[24] = W[24];
  assign P[25] = W[25];
  assign P[26] = W[26];
  assign P[27] = W[27];
  assign P[28] = W[28];
  assign P[29] = W[29];
  MultUB_STD_SD2RBT000 U0 (W, IN1, IN2);
endmodule

module MultUB_STD_SD2RBT000 (P, IN1, IN2);
  output [32:0] P;
  input [14:0] IN1;
  input [14:0] IN2;
  wire [16:0] PP0__dp, PP0__dn;
  wire [18:2] PP1__dp, PP1__dn;
  wire [20:4] PP2__dp, PP2__dn;
  wire [22:6] PP3__dp, PP3__dn;
  wire [24:8] PP4__dp, PP4__dn;
  wire [26:10] PP5__dp, PP5__dn;
  wire [28:12] PP6__dp, PP6__dn;
  wire [28:1] PP7__dp, PP7__dn;
  wire [31:0] Z__dp, Z__dn;
  UBSPPG_14_0_14_0 U0 (PP0__dp, PP0__dn, PP1__dp, PP1__dn, PP2__dp, PP2__dn, PP3__dp, PP3__dn, PP4__dp, PP4__dn, PP5__dp, PP5__dn, PP6__dp, PP6__dn, PP7__dp, PP7__dn, IN1, IN2);
  SD2RBTR_16_0_18_2000 U1 (Z__dp[31:0], Z__dn[31:0], PP0__dp, PP0__dn, PP1__dp, PP1__dn, PP2__dp, PP2__dn, PP3__dp, PP3__dn, PP4__dp, PP4__dn, PP5__dp, PP5__dn, PP6__dp, PP6__dn, PP7__dp, PP7__dn);
  SD2TCConv_FCSkA_3000 U2 (P, Z__dp, Z__dn);
endmodule

module NUBCMBIN_13_13_11000 (O, IN0, IN1, IN2, IN3, IN4, IN5, IN6);
  output [13:1] O;
  input IN0;
  input IN1;
  input IN2;
  input IN3;
  input IN4;
  input IN5;
  input IN6;
  NUB1DCON_13 U0 (O[13], IN0);
  NUBZero_12_12 U1 (O[12]);
  NUB1DCON_11 U2 (O[11], IN1);
  NUBZero_10_10 U3 (O[10]);
  NUB1DCON_9 U4 (O[9], IN2);
  NUBZero_8_8 U5 (O[8]);
  NUB1DCON_7 U6 (O[7], IN3);
  NUBZero_6_6 U7 (O[6]);
  NUB1DCON_5 U8 (O[5], IN4);
  NUBZero_4_4 U9 (O[4]);
  NUB1DCON_3 U10 (O[3], IN5);
  NUBZero_2_2 U11 (O[2]);
  NUB1DCON_1 U12 (O[1], IN6);
endmodule

module NUBCMBIN_16_16_15000 (O, IN0, IN1, IN2);
  output [16:0] O;
  input IN0;
  input [15:1] IN1;
  input IN2;
  NUB1DCON_16 U0 (O[16], IN0);
  NUBCON_15_1 U1 (O[15:1], IN1);
  NUB1DCON_0 U2 (O[0], IN2);
endmodule

module NUBCMBIN_18_18_17000 (O, IN0, IN1, IN2);
  output [18:2] O;
  input IN0;
  input [17:3] IN1;
  input IN2;
  NUB1DCON_18 U0 (O[18], IN0);
  NUBCON_17_3 U1 (O[17:3], IN1);
  NUB1DCON_2 U2 (O[2], IN2);
endmodule

module NUBCMBIN_20_20_19000 (O, IN0, IN1, IN2);
  output [20:4] O;
  input IN0;
  input [19:5] IN1;
  input IN2;
  NUB1DCON_20 U0 (O[20], IN0);
  NUBCON_19_5 U1 (O[19:5], IN1);
  NUB1DCON_4 U2 (O[4], IN2);
endmodule

module NUBCMBIN_22_22_21000 (O, IN0, IN1, IN2);
  output [22:6] O;
  input IN0;
  input [21:7] IN1;
  input IN2;
  NUB1DCON_22 U0 (O[22], IN0);
  NUBCON_21_7 U1 (O[21:7], IN1);
  NUB1DCON_6 U2 (O[6], IN2);
endmodule

module NUBCMBIN_24_24_23000 (O, IN0, IN1, IN2);
  output [24:8] O;
  input IN0;
  input [23:9] IN1;
  input IN2;
  NUB1DCON_24 U0 (O[24], IN0);
  NUBCON_23_9 U1 (O[23:9], IN1);
  NUB1DCON_8 U2 (O[8], IN2);
endmodule

module NUBCMBIN_26_26_25000 (O, IN0, IN1, IN2);
  output [26:10] O;
  input IN0;
  input [25:11] IN1;
  input IN2;
  NUB1DCON_26 U0 (O[26], IN0);
  NUBCON_25_11 U1 (O[25:11], IN1);
  NUB1DCON_10 U2 (O[10], IN2);
endmodule

module NUBCMBIN_28_14_13000 (O, IN0, IN1);
  output [28:1] O;
  input [28:14] IN0;
  input [13:1] IN1;
  NUBCON_28_14 U0 (O[28:14], IN0);
  NUBCON_13_1 U1 (O[13:1], IN1);
endmodule

module NUBCMBIN_28_28_27000 (O, IN0, IN1, IN2);
  output [28:12] O;
  input IN0;
  input [27:13] IN1;
  input IN2;
  NUB1DCON_28 U0 (O[28], IN0);
  NUBCON_27_13 U1 (O[27:13], IN1);
  NUB1DCON_12 U2 (O[12], IN2);
endmodule

module NUBCON_13_1 (O, I);
  output [13:1] O;
  input [13:1] I;
  NUB1DCON_1 U0 (O[1], I[1]);
  NUB1DCON_2 U1 (O[2], I[2]);
  NUB1DCON_3 U2 (O[3], I[3]);
  NUB1DCON_4 U3 (O[4], I[4]);
  NUB1DCON_5 U4 (O[5], I[5]);
  NUB1DCON_6 U5 (O[6], I[6]);
  NUB1DCON_7 U6 (O[7], I[7]);
  NUB1DCON_8 U7 (O[8], I[8]);
  NUB1DCON_9 U8 (O[9], I[9]);
  NUB1DCON_10 U9 (O[10], I[10]);
  NUB1DCON_11 U10 (O[11], I[11]);
  NUB1DCON_12 U11 (O[12], I[12]);
  NUB1DCON_13 U12 (O[13], I[13]);
endmodule

module NUBCON_15_1 (O, I);
  output [15:1] O;
  input [15:1] I;
  NUB1DCON_1 U0 (O[1], I[1]);
  NUB1DCON_2 U1 (O[2], I[2]);
  NUB1DCON_3 U2 (O[3], I[3]);
  NUB1DCON_4 U3 (O[4], I[4]);
  NUB1DCON_5 U4 (O[5], I[5]);
  NUB1DCON_6 U5 (O[6], I[6]);
  NUB1DCON_7 U6 (O[7], I[7]);
  NUB1DCON_8 U7 (O[8], I[8]);
  NUB1DCON_9 U8 (O[9], I[9]);
  NUB1DCON_10 U9 (O[10], I[10]);
  NUB1DCON_11 U10 (O[11], I[11]);
  NUB1DCON_12 U11 (O[12], I[12]);
  NUB1DCON_13 U12 (O[13], I[13]);
  NUB1DCON_14 U13 (O[14], I[14]);
  NUB1DCON_15 U14 (O[15], I[15]);
endmodule

module NUBCON_17_3 (O, I);
  output [17:3] O;
  input [17:3] I;
  NUB1DCON_3 U0 (O[3], I[3]);
  NUB1DCON_4 U1 (O[4], I[4]);
  NUB1DCON_5 U2 (O[5], I[5]);
  NUB1DCON_6 U3 (O[6], I[6]);
  NUB1DCON_7 U4 (O[7], I[7]);
  NUB1DCON_8 U5 (O[8], I[8]);
  NUB1DCON_9 U6 (O[9], I[9]);
  NUB1DCON_10 U7 (O[10], I[10]);
  NUB1DCON_11 U8 (O[11], I[11]);
  NUB1DCON_12 U9 (O[12], I[12]);
  NUB1DCON_13 U10 (O[13], I[13]);
  NUB1DCON_14 U11 (O[14], I[14]);
  NUB1DCON_15 U12 (O[15], I[15]);
  NUB1DCON_16 U13 (O[16], I[16]);
  NUB1DCON_17 U14 (O[17], I[17]);
endmodule

module NUBCON_19_5 (O, I);
  output [19:5] O;
  input [19:5] I;
  NUB1DCON_5 U0 (O[5], I[5]);
  NUB1DCON_6 U1 (O[6], I[6]);
  NUB1DCON_7 U2 (O[7], I[7]);
  NUB1DCON_8 U3 (O[8], I[8]);
  NUB1DCON_9 U4 (O[9], I[9]);
  NUB1DCON_10 U5 (O[10], I[10]);
  NUB1DCON_11 U6 (O[11], I[11]);
  NUB1DCON_12 U7 (O[12], I[12]);
  NUB1DCON_13 U8 (O[13], I[13]);
  NUB1DCON_14 U9 (O[14], I[14]);
  NUB1DCON_15 U10 (O[15], I[15]);
  NUB1DCON_16 U11 (O[16], I[16]);
  NUB1DCON_17 U12 (O[17], I[17]);
  NUB1DCON_18 U13 (O[18], I[18]);
  NUB1DCON_19 U14 (O[19], I[19]);
endmodule

module NUBCON_21_7 (O, I);
  output [21:7] O;
  input [21:7] I;
  NUB1DCON_7 U0 (O[7], I[7]);
  NUB1DCON_8 U1 (O[8], I[8]);
  NUB1DCON_9 U2 (O[9], I[9]);
  NUB1DCON_10 U3 (O[10], I[10]);
  NUB1DCON_11 U4 (O[11], I[11]);
  NUB1DCON_12 U5 (O[12], I[12]);
  NUB1DCON_13 U6 (O[13], I[13]);
  NUB1DCON_14 U7 (O[14], I[14]);
  NUB1DCON_15 U8 (O[15], I[15]);
  NUB1DCON_16 U9 (O[16], I[16]);
  NUB1DCON_17 U10 (O[17], I[17]);
  NUB1DCON_18 U11 (O[18], I[18]);
  NUB1DCON_19 U12 (O[19], I[19]);
  NUB1DCON_20 U13 (O[20], I[20]);
  NUB1DCON_21 U14 (O[21], I[21]);
endmodule

module NUBCON_23_9 (O, I);
  output [23:9] O;
  input [23:9] I;
  NUB1DCON_9 U0 (O[9], I[9]);
  NUB1DCON_10 U1 (O[10], I[10]);
  NUB1DCON_11 U2 (O[11], I[11]);
  NUB1DCON_12 U3 (O[12], I[12]);
  NUB1DCON_13 U4 (O[13], I[13]);
  NUB1DCON_14 U5 (O[14], I[14]);
  NUB1DCON_15 U6 (O[15], I[15]);
  NUB1DCON_16 U7 (O[16], I[16]);
  NUB1DCON_17 U8 (O[17], I[17]);
  NUB1DCON_18 U9 (O[18], I[18]);
  NUB1DCON_19 U10 (O[19], I[19]);
  NUB1DCON_20 U11 (O[20], I[20]);
  NUB1DCON_21 U12 (O[21], I[21]);
  NUB1DCON_22 U13 (O[22], I[22]);
  NUB1DCON_23 U14 (O[23], I[23]);
endmodule

module NUBCON_25_11 (O, I);
  output [25:11] O;
  input [25:11] I;
  NUB1DCON_11 U0 (O[11], I[11]);
  NUB1DCON_12 U1 (O[12], I[12]);
  NUB1DCON_13 U2 (O[13], I[13]);
  NUB1DCON_14 U3 (O[14], I[14]);
  NUB1DCON_15 U4 (O[15], I[15]);
  NUB1DCON_16 U5 (O[16], I[16]);
  NUB1DCON_17 U6 (O[17], I[17]);
  NUB1DCON_18 U7 (O[18], I[18]);
  NUB1DCON_19 U8 (O[19], I[19]);
  NUB1DCON_20 U9 (O[20], I[20]);
  NUB1DCON_21 U10 (O[21], I[21]);
  NUB1DCON_22 U11 (O[22], I[22]);
  NUB1DCON_23 U12 (O[23], I[23]);
  NUB1DCON_24 U13 (O[24], I[24]);
  NUB1DCON_25 U14 (O[25], I[25]);
endmodule

module NUBCON_27_13 (O, I);
  output [27:13] O;
  input [27:13] I;
  NUB1DCON_13 U0 (O[13], I[13]);
  NUB1DCON_14 U1 (O[14], I[14]);
  NUB1DCON_15 U2 (O[15], I[15]);
  NUB1DCON_16 U3 (O[16], I[16]);
  NUB1DCON_17 U4 (O[17], I[17]);
  NUB1DCON_18 U5 (O[18], I[18]);
  NUB1DCON_19 U6 (O[19], I[19]);
  NUB1DCON_20 U7 (O[20], I[20]);
  NUB1DCON_21 U8 (O[21], I[21]);
  NUB1DCON_22 U9 (O[22], I[22]);
  NUB1DCON_23 U10 (O[23], I[23]);
  NUB1DCON_24 U11 (O[24], I[24]);
  NUB1DCON_25 U12 (O[25], I[25]);
  NUB1DCON_26 U13 (O[26], I[26]);
  NUB1DCON_27 U14 (O[27], I[27]);
endmodule

module NUBCON_28_14 (O, I);
  output [28:14] O;
  input [28:14] I;
  NUB1DCON_14 U0 (O[14], I[14]);
  NUB1DCON_15 U1 (O[15], I[15]);
  NUB1DCON_16 U2 (O[16], I[16]);
  NUB1DCON_17 U3 (O[17], I[17]);
  NUB1DCON_18 U4 (O[18], I[18]);
  NUB1DCON_19 U5 (O[19], I[19]);
  NUB1DCON_20 U6 (O[20], I[20]);
  NUB1DCON_21 U7 (O[21], I[21]);
  NUB1DCON_22 U8 (O[22], I[22]);
  NUB1DCON_23 U9 (O[23], I[23]);
  NUB1DCON_24 U10 (O[24], I[24]);
  NUB1DCON_25 U11 (O[25], I[25]);
  NUB1DCON_26 U12 (O[26], I[26]);
  NUB1DCON_27 U13 (O[27], I[27]);
  NUB1DCON_28 U14 (O[28], I[28]);
endmodule

module SD2Decom_PN_31_0 (X, Y, I__dp, I__dn);
  output [31:0] X;
  output [31:0] Y;
  input [31:0] I__dp, I__dn;
  SD2DigitDecom_PN_030 U0 (X[0], Y[0], I__dp[0], I__dn[0]);
  SD2DigitDecom_PN_028 U1 (X[1], Y[1], I__dp[1], I__dn[1]);
  SD2DigitDecom_PN_000 U2 (X[2], Y[2], I__dp[2], I__dn[2]);
  SD2DigitDecom_PN_001 U3 (X[3], Y[3], I__dp[3], I__dn[3]);
  SD2DigitDecom_PN_002 U4 (X[4], Y[4], I__dp[4], I__dn[4]);
  SD2DigitDecom_PN_003 U5 (X[5], Y[5], I__dp[5], I__dn[5]);
  SD2DigitDecom_PN_004 U6 (X[6], Y[6], I__dp[6], I__dn[6]);
  SD2DigitDecom_PN_005 U7 (X[7], Y[7], I__dp[7], I__dn[7]);
  SD2DigitDecom_PN_006 U8 (X[8], Y[8], I__dp[8], I__dn[8]);
  SD2DigitDecom_PN_007 U9 (X[9], Y[9], I__dp[9], I__dn[9]);
  SD2DigitDecom_PN_008 U10 (X[10], Y[10], I__dp[10], I__dn[10]);
  SD2DigitDecom_PN_009 U11 (X[11], Y[11], I__dp[11], I__dn[11]);
  SD2DigitDecom_PN_010 U12 (X[12], Y[12], I__dp[12], I__dn[12]);
  SD2DigitDecom_PN_011 U13 (X[13], Y[13], I__dp[13], I__dn[13]);
  SD2DigitDecom_PN_012 U14 (X[14], Y[14], I__dp[14], I__dn[14]);
  SD2DigitDecom_PN_013 U15 (X[15], Y[15], I__dp[15], I__dn[15]);
  SD2DigitDecom_PN_014 U16 (X[16], Y[16], I__dp[16], I__dn[16]);
  SD2DigitDecom_PN_015 U17 (X[17], Y[17], I__dp[17], I__dn[17]);
  SD2DigitDecom_PN_016 U18 (X[18], Y[18], I__dp[18], I__dn[18]);
  SD2DigitDecom_PN_017 U19 (X[19], Y[19], I__dp[19], I__dn[19]);
  SD2DigitDecom_PN_018 U20 (X[20], Y[20], I__dp[20], I__dn[20]);
  SD2DigitDecom_PN_019 U21 (X[21], Y[21], I__dp[21], I__dn[21]);
  SD2DigitDecom_PN_020 U22 (X[22], Y[22], I__dp[22], I__dn[22]);
  SD2DigitDecom_PN_021 U23 (X[23], Y[23], I__dp[23], I__dn[23]);
  SD2DigitDecom_PN_022 U24 (X[24], Y[24], I__dp[24], I__dn[24]);
  SD2DigitDecom_PN_023 U25 (X[25], Y[25], I__dp[25], I__dn[25]);
  SD2DigitDecom_PN_024 U26 (X[26], Y[26], I__dp[26], I__dn[26]);
  SD2DigitDecom_PN_025 U27 (X[27], Y[27], I__dp[27], I__dn[27]);
  SD2DigitDecom_PN_026 U28 (X[28], Y[28], I__dp[28], I__dn[28]);
  SD2DigitDecom_PN_027 U29 (X[29], Y[29], I__dp[29], I__dn[29]);
  SD2DigitDecom_PN_029 U30 (X[30], Y[30], I__dp[30], I__dn[30]);
  SD2DigitDecom_PN_031 U31 (X[31], Y[31], I__dp[31], I__dn[31]);
endmodule

module SD2DigitRBA_1 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_028 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_028 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_1 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_1 U3 (C2, S2, C1i, S1, Yp);
  UBInv_2 U4 (C2o, C2);
  SD2DigitCom_1 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_10 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_008 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_008 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_10 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_10 U3 (C2, S2, C1i, S1, Yp);
  UBInv_11 U4 (C2o, C2);
  SD2DigitCom_10 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_11 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_009 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_009 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_11 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_11 U3 (C2, S2, C1i, S1, Yp);
  UBInv_12 U4 (C2o, C2);
  SD2DigitCom_11 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_12 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_010 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_010 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_12 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_12 U3 (C2, S2, C1i, S1, Yp);
  UBInv_13 U4 (C2o, C2);
  SD2DigitCom_12 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_13 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_011 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_011 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_13 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_13 U3 (C2, S2, C1i, S1, Yp);
  UBInv_14 U4 (C2o, C2);
  SD2DigitCom_13 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_14 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_012 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_012 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_14 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_14 U3 (C2, S2, C1i, S1, Yp);
  UBInv_15 U4 (C2o, C2);
  SD2DigitCom_14 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_15 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_013 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_013 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_15 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_15 U3 (C2, S2, C1i, S1, Yp);
  UBInv_16 U4 (C2o, C2);
  SD2DigitCom_15 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_16 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_014 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_014 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_16 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_16 U3 (C2, S2, C1i, S1, Yp);
  UBInv_17 U4 (C2o, C2);
  SD2DigitCom_16 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_17 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_015 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_015 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_17 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_17 U3 (C2, S2, C1i, S1, Yp);
  UBInv_18 U4 (C2o, C2);
  SD2DigitCom_17 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_18 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_016 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_016 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_18 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_18 U3 (C2, S2, C1i, S1, Yp);
  UBInv_19 U4 (C2o, C2);
  SD2DigitCom_18 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_19 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_017 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_017 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_19 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_19 U3 (C2, S2, C1i, S1, Yp);
  UBInv_20 U4 (C2o, C2);
  SD2DigitCom_19 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_2 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_000 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_000 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_2 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_2 U3 (C2, S2, C1i, S1, Yp);
  UBInv_3 U4 (C2o, C2);
  SD2DigitCom_2 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_20 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_018 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_018 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_20 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_20 U3 (C2, S2, C1i, S1, Yp);
  UBInv_21 U4 (C2o, C2);
  SD2DigitCom_20 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_21 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_019 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_019 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_21 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_21 U3 (C2, S2, C1i, S1, Yp);
  UBInv_22 U4 (C2o, C2);
  SD2DigitCom_21 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_22 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_020 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_020 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_22 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_22 U3 (C2, S2, C1i, S1, Yp);
  UBInv_23 U4 (C2o, C2);
  SD2DigitCom_22 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_23 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_021 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_021 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_23 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_23 U3 (C2, S2, C1i, S1, Yp);
  UBInv_24 U4 (C2o, C2);
  SD2DigitCom_23 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_24 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_022 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_022 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_24 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_24 U3 (C2, S2, C1i, S1, Yp);
  UBInv_25 U4 (C2o, C2);
  SD2DigitCom_24 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_25 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_023 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_023 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_25 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_25 U3 (C2, S2, C1i, S1, Yp);
  UBInv_26 U4 (C2o, C2);
  SD2DigitCom_25 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_26 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_024 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_024 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_26 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_26 U3 (C2, S2, C1i, S1, Yp);
  UBInv_27 U4 (C2o, C2);
  SD2DigitCom_26 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_27 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_025 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_025 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_27 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_27 U3 (C2, S2, C1i, S1, Yp);
  UBInv_28 U4 (C2o, C2);
  SD2DigitCom_27 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_28 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_026 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_026 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_28 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_28 U3 (C2, S2, C1i, S1, Yp);
  UBInv_29 U4 (C2o, C2);
  SD2DigitCom_28 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_29 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_027 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_027 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_29 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_29 U3 (C2, S2, C1i, S1, Yp);
  UBInv_30 U4 (C2o, C2);
  SD2DigitCom_29 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_3 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_001 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_001 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_3 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_3 U3 (C2, S2, C1i, S1, Yp);
  UBInv_4 U4 (C2o, C2);
  SD2DigitCom_3 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_30 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_029 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_029 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_30 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_30 U3 (C2, S2, C1i, S1, Yp);
  UBInv_31 U4 (C2o, C2);
  SD2DigitCom_30 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_4 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_002 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_002 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_4 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_4 U3 (C2, S2, C1i, S1, Yp);
  UBInv_5 U4 (C2o, C2);
  SD2DigitCom_4 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_5 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_003 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_003 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_5 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_5 U3 (C2, S2, C1i, S1, Yp);
  UBInv_6 U4 (C2o, C2);
  SD2DigitCom_5 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_6 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_004 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_004 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_6 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_6 U3 (C2, S2, C1i, S1, Yp);
  UBInv_7 U4 (C2o, C2);
  SD2DigitCom_6 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_7 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_005 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_005 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_7 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_7 U3 (C2, S2, C1i, S1, Yp);
  UBInv_8 U4 (C2o, C2);
  SD2DigitCom_7 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_8 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_006 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_006 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_8 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_8 U3 (C2, S2, C1i, S1, Yp);
  UBInv_9 U4 (C2o, C2);
  SD2DigitCom_8 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2DigitRBA_9 (Z__dp, Z__dn, C1o, C2o, X__dp, X__dn, Y__dp, Y__dn, C1i, C2i);
  output C1o;
  output C2o;
  output Z__dp, Z__dn;
  input C1i;
  input C2i;
  input X__dp, X__dn;
  input Y__dp, Y__dn;
  wire C2;
  wire S1;
  wire S2;
  wire Xn;
  wire Xp;
  wire Yn;
  wire Yp;
  SD2DigitDecom_PN_007 U0 (Xn, Xp, X__dp, X__dn);
  SD2DigitDecom_PN_007 U1 (Yn, Yp, Y__dp, Y__dn);
  UBFA_9 U2 (C1o, S1, Xn, Xp, Yn);
  UBFA_9 U3 (C2, S2, C1i, S1, Yp);
  UBInv_10 U4 (C2o, C2);
  SD2DigitCom_9 U5 (Z__dp, Z__dn, C2i, S2);
endmodule

module SD2PureRBA_18_2 (Z__dp, Z__dn, X__dp, X__dn, Y__dp, Y__dn);
  output [19:2] Z__dp, Z__dn;
  input [18:2] X__dp, X__dn;
  input [18:2] Y__dp, Y__dn;
  wire C1_10;
  wire C1_11;
  wire C1_12;
  wire C1_13;
  wire C1_14;
  wire C1_15;
  wire C1_16;
  wire C1_17;
  wire C1_18;
  wire C1_19;
  wire C1_3;
  wire C1_4;
  wire C1_5;
  wire C1_6;
  wire C1_7;
  wire C1_8;
  wire C1_9;
  wire C1i;
  wire C2_10;
  wire C2_11;
  wire C2_12;
  wire C2_13;
  wire C2_14;
  wire C2_15;
  wire C2_16;
  wire C2_17;
  wire C2_18;
  wire C2_19;
  wire C2_3;
  wire C2_4;
  wire C2_5;
  wire C2_6;
  wire C2_7;
  wire C2_8;
  wire C2_9;
  wire C2i;
  UBZero_2_2 U0 (C1i);
  NUBZero_2_2 U1 (C2i);
  SD2DigitRBA_2 U2 (Z__dp[2], Z__dn[2], C1_3, C2_3, X__dp[2], X__dn[2], Y__dp[2], Y__dn[2], C1i, C2i);
  SD2DigitRBA_3 U3 (Z__dp[3], Z__dn[3], C1_4, C2_4, X__dp[3], X__dn[3], Y__dp[3], Y__dn[3], C1_3, C2_3);
  SD2DigitRBA_4 U4 (Z__dp[4], Z__dn[4], C1_5, C2_5, X__dp[4], X__dn[4], Y__dp[4], Y__dn[4], C1_4, C2_4);
  SD2DigitRBA_5 U5 (Z__dp[5], Z__dn[5], C1_6, C2_6, X__dp[5], X__dn[5], Y__dp[5], Y__dn[5], C1_5, C2_5);
  SD2DigitRBA_6 U6 (Z__dp[6], Z__dn[6], C1_7, C2_7, X__dp[6], X__dn[6], Y__dp[6], Y__dn[6], C1_6, C2_6);
  SD2DigitRBA_7 U7 (Z__dp[7], Z__dn[7], C1_8, C2_8, X__dp[7], X__dn[7], Y__dp[7], Y__dn[7], C1_7, C2_7);
  SD2DigitRBA_8 U8 (Z__dp[8], Z__dn[8], C1_9, C2_9, X__dp[8], X__dn[8], Y__dp[8], Y__dn[8], C1_8, C2_8);
  SD2DigitRBA_9 U9 (Z__dp[9], Z__dn[9], C1_10, C2_10, X__dp[9], X__dn[9], Y__dp[9], Y__dn[9], C1_9, C2_9);
  SD2DigitRBA_10 U10 (Z__dp[10], Z__dn[10], C1_11, C2_11, X__dp[10], X__dn[10], Y__dp[10], Y__dn[10], C1_10, C2_10);
  SD2DigitRBA_11 U11 (Z__dp[11], Z__dn[11], C1_12, C2_12, X__dp[11], X__dn[11], Y__dp[11], Y__dn[11], C1_11, C2_11);
  SD2DigitRBA_12 U12 (Z__dp[12], Z__dn[12], C1_13, C2_13, X__dp[12], X__dn[12], Y__dp[12], Y__dn[12], C1_12, C2_12);
  SD2DigitRBA_13 U13 (Z__dp[13], Z__dn[13], C1_14, C2_14, X__dp[13], X__dn[13], Y__dp[13], Y__dn[13], C1_13, C2_13);
  SD2DigitRBA_14 U14 (Z__dp[14], Z__dn[14], C1_15, C2_15, X__dp[14], X__dn[14], Y__dp[14], Y__dn[14], C1_14, C2_14);
  SD2DigitRBA_15 U15 (Z__dp[15], Z__dn[15], C1_16, C2_16, X__dp[15], X__dn[15], Y__dp[15], Y__dn[15], C1_15, C2_15);
  SD2DigitRBA_16 U16 (Z__dp[16], Z__dn[16], C1_17, C2_17, X__dp[16], X__dn[16], Y__dp[16], Y__dn[16], C1_16, C2_16);
  SD2DigitRBA_17 U17 (Z__dp[17], Z__dn[17], C1_18, C2_18, X__dp[17], X__dn[17], Y__dp[17], Y__dn[17], C1_17, C2_17);
  SD2DigitRBA_18 U18 (Z__dp[18], Z__dn[18], C1_19, C2_19, X__dp[18], X__dn[18], Y__dp[18], Y__dn[18], C1_18, C2_18);
  SD2DigitCom_19 U19 (Z__dp[19], Z__dn[19], C2_19, C1_19);
endmodule

module SD2PureRBA_22_6 (Z__dp, Z__dn, X__dp, X__dn, Y__dp, Y__dn);
  output [23:6] Z__dp, Z__dn;
  input [22:6] X__dp, X__dn;
  input [22:6] Y__dp, Y__dn;
  wire C1_10;
  wire C1_11;
  wire C1_12;
  wire C1_13;
  wire C1_14;
  wire C1_15;
  wire C1_16;
  wire C1_17;
  wire C1_18;
  wire C1_19;
  wire C1_20;
  wire C1_21;
  wire C1_22;
  wire C1_23;
  wire C1_7;
  wire C1_8;
  wire C1_9;
  wire C1i;
  wire C2_10;
  wire C2_11;
  wire C2_12;
  wire C2_13;
  wire C2_14;
  wire C2_15;
  wire C2_16;
  wire C2_17;
  wire C2_18;
  wire C2_19;
  wire C2_20;
  wire C2_21;
  wire C2_22;
  wire C2_23;
  wire C2_7;
  wire C2_8;
  wire C2_9;
  wire C2i;
  UBZero_6_6 U0 (C1i);
  NUBZero_6_6 U1 (C2i);
  SD2DigitRBA_6 U2 (Z__dp[6], Z__dn[6], C1_7, C2_7, X__dp[6], X__dn[6], Y__dp[6], Y__dn[6], C1i, C2i);
  SD2DigitRBA_7 U3 (Z__dp[7], Z__dn[7], C1_8, C2_8, X__dp[7], X__dn[7], Y__dp[7], Y__dn[7], C1_7, C2_7);
  SD2DigitRBA_8 U4 (Z__dp[8], Z__dn[8], C1_9, C2_9, X__dp[8], X__dn[8], Y__dp[8], Y__dn[8], C1_8, C2_8);
  SD2DigitRBA_9 U5 (Z__dp[9], Z__dn[9], C1_10, C2_10, X__dp[9], X__dn[9], Y__dp[9], Y__dn[9], C1_9, C2_9);
  SD2DigitRBA_10 U6 (Z__dp[10], Z__dn[10], C1_11, C2_11, X__dp[10], X__dn[10], Y__dp[10], Y__dn[10], C1_10, C2_10);
  SD2DigitRBA_11 U7 (Z__dp[11], Z__dn[11], C1_12, C2_12, X__dp[11], X__dn[11], Y__dp[11], Y__dn[11], C1_11, C2_11);
  SD2DigitRBA_12 U8 (Z__dp[12], Z__dn[12], C1_13, C2_13, X__dp[12], X__dn[12], Y__dp[12], Y__dn[12], C1_12, C2_12);
  SD2DigitRBA_13 U9 (Z__dp[13], Z__dn[13], C1_14, C2_14, X__dp[13], X__dn[13], Y__dp[13], Y__dn[13], C1_13, C2_13);
  SD2DigitRBA_14 U10 (Z__dp[14], Z__dn[14], C1_15, C2_15, X__dp[14], X__dn[14], Y__dp[14], Y__dn[14], C1_14, C2_14);
  SD2DigitRBA_15 U11 (Z__dp[15], Z__dn[15], C1_16, C2_16, X__dp[15], X__dn[15], Y__dp[15], Y__dn[15], C1_15, C2_15);
  SD2DigitRBA_16 U12 (Z__dp[16], Z__dn[16], C1_17, C2_17, X__dp[16], X__dn[16], Y__dp[16], Y__dn[16], C1_16, C2_16);
  SD2DigitRBA_17 U13 (Z__dp[17], Z__dn[17], C1_18, C2_18, X__dp[17], X__dn[17], Y__dp[17], Y__dn[17], C1_17, C2_17);
  SD2DigitRBA_18 U14 (Z__dp[18], Z__dn[18], C1_19, C2_19, X__dp[18], X__dn[18], Y__dp[18], Y__dn[18], C1_18, C2_18);
  SD2DigitRBA_19 U15 (Z__dp[19], Z__dn[19], C1_20, C2_20, X__dp[19], X__dn[19], Y__dp[19], Y__dn[19], C1_19, C2_19);
  SD2DigitRBA_20 U16 (Z__dp[20], Z__dn[20], C1_21, C2_21, X__dp[20], X__dn[20], Y__dp[20], Y__dn[20], C1_20, C2_20);
  SD2DigitRBA_21 U17 (Z__dp[21], Z__dn[21], C1_22, C2_22, X__dp[21], X__dn[21], Y__dp[21], Y__dn[21], C1_21, C2_21);
  SD2DigitRBA_22 U18 (Z__dp[22], Z__dn[22], C1_23, C2_23, X__dp[22], X__dn[22], Y__dp[22], Y__dn[22], C1_22, C2_22);
  SD2DigitCom_23 U19 (Z__dp[23], Z__dn[23], C2_23, C1_23);
endmodule

module SD2PureRBA_23_4 (Z__dp, Z__dn, X__dp, X__dn, Y__dp, Y__dn);
  output [24:4] Z__dp, Z__dn;
  input [23:4] X__dp, X__dn;
  input [23:4] Y__dp, Y__dn;
  wire C1_10;
  wire C1_11;
  wire C1_12;
  wire C1_13;
  wire C1_14;
  wire C1_15;
  wire C1_16;
  wire C1_17;
  wire C1_18;
  wire C1_19;
  wire C1_20;
  wire C1_21;
  wire C1_22;
  wire C1_23;
  wire C1_24;
  wire C1_5;
  wire C1_6;
  wire C1_7;
  wire C1_8;
  wire C1_9;
  wire C1i;
  wire C2_10;
  wire C2_11;
  wire C2_12;
  wire C2_13;
  wire C2_14;
  wire C2_15;
  wire C2_16;
  wire C2_17;
  wire C2_18;
  wire C2_19;
  wire C2_20;
  wire C2_21;
  wire C2_22;
  wire C2_23;
  wire C2_24;
  wire C2_5;
  wire C2_6;
  wire C2_7;
  wire C2_8;
  wire C2_9;
  wire C2i;
  UBZero_4_4 U0 (C1i);
  NUBZero_4_4 U1 (C2i);
  SD2DigitRBA_4 U2 (Z__dp[4], Z__dn[4], C1_5, C2_5, X__dp[4], X__dn[4], Y__dp[4], Y__dn[4], C1i, C2i);
  SD2DigitRBA_5 U3 (Z__dp[5], Z__dn[5], C1_6, C2_6, X__dp[5], X__dn[5], Y__dp[5], Y__dn[5], C1_5, C2_5);
  SD2DigitRBA_6 U4 (Z__dp[6], Z__dn[6], C1_7, C2_7, X__dp[6], X__dn[6], Y__dp[6], Y__dn[6], C1_6, C2_6);
  SD2DigitRBA_7 U5 (Z__dp[7], Z__dn[7], C1_8, C2_8, X__dp[7], X__dn[7], Y__dp[7], Y__dn[7], C1_7, C2_7);
  SD2DigitRBA_8 U6 (Z__dp[8], Z__dn[8], C1_9, C2_9, X__dp[8], X__dn[8], Y__dp[8], Y__dn[8], C1_8, C2_8);
  SD2DigitRBA_9 U7 (Z__dp[9], Z__dn[9], C1_10, C2_10, X__dp[9], X__dn[9], Y__dp[9], Y__dn[9], C1_9, C2_9);
  SD2DigitRBA_10 U8 (Z__dp[10], Z__dn[10], C1_11, C2_11, X__dp[10], X__dn[10], Y__dp[10], Y__dn[10], C1_10, C2_10);
  SD2DigitRBA_11 U9 (Z__dp[11], Z__dn[11], C1_12, C2_12, X__dp[11], X__dn[11], Y__dp[11], Y__dn[11], C1_11, C2_11);
  SD2DigitRBA_12 U10 (Z__dp[12], Z__dn[12], C1_13, C2_13, X__dp[12], X__dn[12], Y__dp[12], Y__dn[12], C1_12, C2_12);
  SD2DigitRBA_13 U11 (Z__dp[13], Z__dn[13], C1_14, C2_14, X__dp[13], X__dn[13], Y__dp[13], Y__dn[13], C1_13, C2_13);
  SD2DigitRBA_14 U12 (Z__dp[14], Z__dn[14], C1_15, C2_15, X__dp[14], X__dn[14], Y__dp[14], Y__dn[14], C1_14, C2_14);
  SD2DigitRBA_15 U13 (Z__dp[15], Z__dn[15], C1_16, C2_16, X__dp[15], X__dn[15], Y__dp[15], Y__dn[15], C1_15, C2_15);
  SD2DigitRBA_16 U14 (Z__dp[16], Z__dn[16], C1_17, C2_17, X__dp[16], X__dn[16], Y__dp[16], Y__dn[16], C1_16, C2_16);
  SD2DigitRBA_17 U15 (Z__dp[17], Z__dn[17], C1_18, C2_18, X__dp[17], X__dn[17], Y__dp[17], Y__dn[17], C1_17, C2_17);
  SD2DigitRBA_18 U16 (Z__dp[18], Z__dn[18], C1_19, C2_19, X__dp[18], X__dn[18], Y__dp[18], Y__dn[18], C1_18, C2_18);
  SD2DigitRBA_19 U17 (Z__dp[19], Z__dn[19], C1_20, C2_20, X__dp[19], X__dn[19], Y__dp[19], Y__dn[19], C1_19, C2_19);
  SD2DigitRBA_20 U18 (Z__dp[20], Z__dn[20], C1_21, C2_21, X__dp[20], X__dn[20], Y__dp[20], Y__dn[20], C1_20, C2_20);
  SD2DigitRBA_21 U19 (Z__dp[21], Z__dn[21], C1_22, C2_22, X__dp[21], X__dn[21], Y__dp[21], Y__dn[21], C1_21, C2_21);
  SD2DigitRBA_22 U20 (Z__dp[22], Z__dn[22], C1_23, C2_23, X__dp[22], X__dn[22], Y__dp[22], Y__dn[22], C1_22, C2_22);
  SD2DigitRBA_23 U21 (Z__dp[23], Z__dn[23], C1_24, C2_24, X__dp[23], X__dn[23], Y__dp[23], Y__dn[23], C1_23, C2_23);
  SD2DigitCom_24 U22 (Z__dp[24], Z__dn[24], C2_24, C1_24);
endmodule

module SD2PureRBA_26_10 (Z__dp, Z__dn, X__dp, X__dn, Y__dp, Y__dn);
  output [27:10] Z__dp, Z__dn;
  input [26:10] X__dp, X__dn;
  input [26:10] Y__dp, Y__dn;
  wire C1_11;
  wire C1_12;
  wire C1_13;
  wire C1_14;
  wire C1_15;
  wire C1_16;
  wire C1_17;
  wire C1_18;
  wire C1_19;
  wire C1_20;
  wire C1_21;
  wire C1_22;
  wire C1_23;
  wire C1_24;
  wire C1_25;
  wire C1_26;
  wire C1_27;
  wire C1i;
  wire C2_11;
  wire C2_12;
  wire C2_13;
  wire C2_14;
  wire C2_15;
  wire C2_16;
  wire C2_17;
  wire C2_18;
  wire C2_19;
  wire C2_20;
  wire C2_21;
  wire C2_22;
  wire C2_23;
  wire C2_24;
  wire C2_25;
  wire C2_26;
  wire C2_27;
  wire C2i;
  UBZero_10_10 U0 (C1i);
  NUBZero_10_10 U1 (C2i);
  SD2DigitRBA_10 U2 (Z__dp[10], Z__dn[10], C1_11, C2_11, X__dp[10], X__dn[10], Y__dp[10], Y__dn[10], C1i, C2i);
  SD2DigitRBA_11 U3 (Z__dp[11], Z__dn[11], C1_12, C2_12, X__dp[11], X__dn[11], Y__dp[11], Y__dn[11], C1_11, C2_11);
  SD2DigitRBA_12 U4 (Z__dp[12], Z__dn[12], C1_13, C2_13, X__dp[12], X__dn[12], Y__dp[12], Y__dn[12], C1_12, C2_12);
  SD2DigitRBA_13 U5 (Z__dp[13], Z__dn[13], C1_14, C2_14, X__dp[13], X__dn[13], Y__dp[13], Y__dn[13], C1_13, C2_13);
  SD2DigitRBA_14 U6 (Z__dp[14], Z__dn[14], C1_15, C2_15, X__dp[14], X__dn[14], Y__dp[14], Y__dn[14], C1_14, C2_14);
  SD2DigitRBA_15 U7 (Z__dp[15], Z__dn[15], C1_16, C2_16, X__dp[15], X__dn[15], Y__dp[15], Y__dn[15], C1_15, C2_15);
  SD2DigitRBA_16 U8 (Z__dp[16], Z__dn[16], C1_17, C2_17, X__dp[16], X__dn[16], Y__dp[16], Y__dn[16], C1_16, C2_16);
  SD2DigitRBA_17 U9 (Z__dp[17], Z__dn[17], C1_18, C2_18, X__dp[17], X__dn[17], Y__dp[17], Y__dn[17], C1_17, C2_17);
  SD2DigitRBA_18 U10 (Z__dp[18], Z__dn[18], C1_19, C2_19, X__dp[18], X__dn[18], Y__dp[18], Y__dn[18], C1_18, C2_18);
  SD2DigitRBA_19 U11 (Z__dp[19], Z__dn[19], C1_20, C2_20, X__dp[19], X__dn[19], Y__dp[19], Y__dn[19], C1_19, C2_19);
  SD2DigitRBA_20 U12 (Z__dp[20], Z__dn[20], C1_21, C2_21, X__dp[20], X__dn[20], Y__dp[20], Y__dn[20], C1_20, C2_20);
  SD2DigitRBA_21 U13 (Z__dp[21], Z__dn[21], C1_22, C2_22, X__dp[21], X__dn[21], Y__dp[21], Y__dn[21], C1_21, C2_21);
  SD2DigitRBA_22 U14 (Z__dp[22], Z__dn[22], C1_23, C2_23, X__dp[22], X__dn[22], Y__dp[22], Y__dn[22], C1_22, C2_22);
  SD2DigitRBA_23 U15 (Z__dp[23], Z__dn[23], C1_24, C2_24, X__dp[23], X__dn[23], Y__dp[23], Y__dn[23], C1_23, C2_23);
  SD2DigitRBA_24 U16 (Z__dp[24], Z__dn[24], C1_25, C2_25, X__dp[24], X__dn[24], Y__dp[24], Y__dn[24], C1_24, C2_24);
  SD2DigitRBA_25 U17 (Z__dp[25], Z__dn[25], C1_26, C2_26, X__dp[25], X__dn[25], Y__dp[25], Y__dn[25], C1_25, C2_25);
  SD2DigitRBA_26 U18 (Z__dp[26], Z__dn[26], C1_27, C2_27, X__dp[26], X__dn[26], Y__dp[26], Y__dn[26], C1_26, C2_26);
  SD2DigitCom_27 U19 (Z__dp[27], Z__dn[27], C2_27, C1_27);
endmodule

module SD2PureRBA_28_12 (Z__dp, Z__dn, X__dp, X__dn, Y__dp, Y__dn);
  output [29:12] Z__dp, Z__dn;
  input [28:12] X__dp, X__dn;
  input [28:12] Y__dp, Y__dn;
  wire C1_13;
  wire C1_14;
  wire C1_15;
  wire C1_16;
  wire C1_17;
  wire C1_18;
  wire C1_19;
  wire C1_20;
  wire C1_21;
  wire C1_22;
  wire C1_23;
  wire C1_24;
  wire C1_25;
  wire C1_26;
  wire C1_27;
  wire C1_28;
  wire C1_29;
  wire C1i;
  wire C2_13;
  wire C2_14;
  wire C2_15;
  wire C2_16;
  wire C2_17;
  wire C2_18;
  wire C2_19;
  wire C2_20;
  wire C2_21;
  wire C2_22;
  wire C2_23;
  wire C2_24;
  wire C2_25;
  wire C2_26;
  wire C2_27;
  wire C2_28;
  wire C2_29;
  wire C2i;
  UBZero_12_12 U0 (C1i);
  NUBZero_12_12 U1 (C2i);
  SD2DigitRBA_12 U2 (Z__dp[12], Z__dn[12], C1_13, C2_13, X__dp[12], X__dn[12], Y__dp[12], Y__dn[12], C1i, C2i);
  SD2DigitRBA_13 U3 (Z__dp[13], Z__dn[13], C1_14, C2_14, X__dp[13], X__dn[13], Y__dp[13], Y__dn[13], C1_13, C2_13);
  SD2DigitRBA_14 U4 (Z__dp[14], Z__dn[14], C1_15, C2_15, X__dp[14], X__dn[14], Y__dp[14], Y__dn[14], C1_14, C2_14);
  SD2DigitRBA_15 U5 (Z__dp[15], Z__dn[15], C1_16, C2_16, X__dp[15], X__dn[15], Y__dp[15], Y__dn[15], C1_15, C2_15);
  SD2DigitRBA_16 U6 (Z__dp[16], Z__dn[16], C1_17, C2_17, X__dp[16], X__dn[16], Y__dp[16], Y__dn[16], C1_16, C2_16);
  SD2DigitRBA_17 U7 (Z__dp[17], Z__dn[17], C1_18, C2_18, X__dp[17], X__dn[17], Y__dp[17], Y__dn[17], C1_17, C2_17);
  SD2DigitRBA_18 U8 (Z__dp[18], Z__dn[18], C1_19, C2_19, X__dp[18], X__dn[18], Y__dp[18], Y__dn[18], C1_18, C2_18);
  SD2DigitRBA_19 U9 (Z__dp[19], Z__dn[19], C1_20, C2_20, X__dp[19], X__dn[19], Y__dp[19], Y__dn[19], C1_19, C2_19);
  SD2DigitRBA_20 U10 (Z__dp[20], Z__dn[20], C1_21, C2_21, X__dp[20], X__dn[20], Y__dp[20], Y__dn[20], C1_20, C2_20);
  SD2DigitRBA_21 U11 (Z__dp[21], Z__dn[21], C1_22, C2_22, X__dp[21], X__dn[21], Y__dp[21], Y__dn[21], C1_21, C2_21);
  SD2DigitRBA_22 U12 (Z__dp[22], Z__dn[22], C1_23, C2_23, X__dp[22], X__dn[22], Y__dp[22], Y__dn[22], C1_22, C2_22);
  SD2DigitRBA_23 U13 (Z__dp[23], Z__dn[23], C1_24, C2_24, X__dp[23], X__dn[23], Y__dp[23], Y__dn[23], C1_23, C2_23);
  SD2DigitRBA_24 U14 (Z__dp[24], Z__dn[24], C1_25, C2_25, X__dp[24], X__dn[24], Y__dp[24], Y__dn[24], C1_24, C2_24);
  SD2DigitRBA_25 U15 (Z__dp[25], Z__dn[25], C1_26, C2_26, X__dp[25], X__dn[25], Y__dp[25], Y__dn[25], C1_25, C2_25);
  SD2DigitRBA_26 U16 (Z__dp[26], Z__dn[26], C1_27, C2_27, X__dp[26], X__dn[26], Y__dp[26], Y__dn[26], C1_26, C2_26);
  SD2DigitRBA_27 U17 (Z__dp[27], Z__dn[27], C1_28, C2_28, X__dp[27], X__dn[27], Y__dp[27], Y__dn[27], C1_27, C2_27);
  SD2DigitRBA_28 U18 (Z__dp[28], Z__dn[28], C1_29, C2_29, X__dp[28], X__dn[28], Y__dp[28], Y__dn[28], C1_28, C2_28);
  SD2DigitCom_29 U19 (Z__dp[29], Z__dn[29], C2_29, C1_29);
endmodule

module SD2PureRBA_29_8 (Z__dp, Z__dn, X__dp, X__dn, Y__dp, Y__dn);
  output [30:8] Z__dp, Z__dn;
  input [29:8] X__dp, X__dn;
  input [29:8] Y__dp, Y__dn;
  wire C1_10;
  wire C1_11;
  wire C1_12;
  wire C1_13;
  wire C1_14;
  wire C1_15;
  wire C1_16;
  wire C1_17;
  wire C1_18;
  wire C1_19;
  wire C1_20;
  wire C1_21;
  wire C1_22;
  wire C1_23;
  wire C1_24;
  wire C1_25;
  wire C1_26;
  wire C1_27;
  wire C1_28;
  wire C1_29;
  wire C1_30;
  wire C1_9;
  wire C1i;
  wire C2_10;
  wire C2_11;
  wire C2_12;
  wire C2_13;
  wire C2_14;
  wire C2_15;
  wire C2_16;
  wire C2_17;
  wire C2_18;
  wire C2_19;
  wire C2_20;
  wire C2_21;
  wire C2_22;
  wire C2_23;
  wire C2_24;
  wire C2_25;
  wire C2_26;
  wire C2_27;
  wire C2_28;
  wire C2_29;
  wire C2_30;
  wire C2_9;
  wire C2i;
  UBZero_8_8 U0 (C1i);
  NUBZero_8_8 U1 (C2i);
  SD2DigitRBA_8 U2 (Z__dp[8], Z__dn[8], C1_9, C2_9, X__dp[8], X__dn[8], Y__dp[8], Y__dn[8], C1i, C2i);
  SD2DigitRBA_9 U3 (Z__dp[9], Z__dn[9], C1_10, C2_10, X__dp[9], X__dn[9], Y__dp[9], Y__dn[9], C1_9, C2_9);
  SD2DigitRBA_10 U4 (Z__dp[10], Z__dn[10], C1_11, C2_11, X__dp[10], X__dn[10], Y__dp[10], Y__dn[10], C1_10, C2_10);
  SD2DigitRBA_11 U5 (Z__dp[11], Z__dn[11], C1_12, C2_12, X__dp[11], X__dn[11], Y__dp[11], Y__dn[11], C1_11, C2_11);
  SD2DigitRBA_12 U6 (Z__dp[12], Z__dn[12], C1_13, C2_13, X__dp[12], X__dn[12], Y__dp[12], Y__dn[12], C1_12, C2_12);
  SD2DigitRBA_13 U7 (Z__dp[13], Z__dn[13], C1_14, C2_14, X__dp[13], X__dn[13], Y__dp[13], Y__dn[13], C1_13, C2_13);
  SD2DigitRBA_14 U8 (Z__dp[14], Z__dn[14], C1_15, C2_15, X__dp[14], X__dn[14], Y__dp[14], Y__dn[14], C1_14, C2_14);
  SD2DigitRBA_15 U9 (Z__dp[15], Z__dn[15], C1_16, C2_16, X__dp[15], X__dn[15], Y__dp[15], Y__dn[15], C1_15, C2_15);
  SD2DigitRBA_16 U10 (Z__dp[16], Z__dn[16], C1_17, C2_17, X__dp[16], X__dn[16], Y__dp[16], Y__dn[16], C1_16, C2_16);
  SD2DigitRBA_17 U11 (Z__dp[17], Z__dn[17], C1_18, C2_18, X__dp[17], X__dn[17], Y__dp[17], Y__dn[17], C1_17, C2_17);
  SD2DigitRBA_18 U12 (Z__dp[18], Z__dn[18], C1_19, C2_19, X__dp[18], X__dn[18], Y__dp[18], Y__dn[18], C1_18, C2_18);
  SD2DigitRBA_19 U13 (Z__dp[19], Z__dn[19], C1_20, C2_20, X__dp[19], X__dn[19], Y__dp[19], Y__dn[19], C1_19, C2_19);
  SD2DigitRBA_20 U14 (Z__dp[20], Z__dn[20], C1_21, C2_21, X__dp[20], X__dn[20], Y__dp[20], Y__dn[20], C1_20, C2_20);
  SD2DigitRBA_21 U15 (Z__dp[21], Z__dn[21], C1_22, C2_22, X__dp[21], X__dn[21], Y__dp[21], Y__dn[21], C1_21, C2_21);
  SD2DigitRBA_22 U16 (Z__dp[22], Z__dn[22], C1_23, C2_23, X__dp[22], X__dn[22], Y__dp[22], Y__dn[22], C1_22, C2_22);
  SD2DigitRBA_23 U17 (Z__dp[23], Z__dn[23], C1_24, C2_24, X__dp[23], X__dn[23], Y__dp[23], Y__dn[23], C1_23, C2_23);
  SD2DigitRBA_24 U18 (Z__dp[24], Z__dn[24], C1_25, C2_25, X__dp[24], X__dn[24], Y__dp[24], Y__dn[24], C1_24, C2_24);
  SD2DigitRBA_25 U19 (Z__dp[25], Z__dn[25], C1_26, C2_26, X__dp[25], X__dn[25], Y__dp[25], Y__dn[25], C1_25, C2_25);
  SD2DigitRBA_26 U20 (Z__dp[26], Z__dn[26], C1_27, C2_27, X__dp[26], X__dn[26], Y__dp[26], Y__dn[26], C1_26, C2_26);
  SD2DigitRBA_27 U21 (Z__dp[27], Z__dn[27], C1_28, C2_28, X__dp[27], X__dn[27], Y__dp[27], Y__dn[27], C1_27, C2_27);
  SD2DigitRBA_28 U22 (Z__dp[28], Z__dn[28], C1_29, C2_29, X__dp[28], X__dn[28], Y__dp[28], Y__dn[28], C1_28, C2_28);
  SD2DigitRBA_29 U23 (Z__dp[29], Z__dn[29], C1_30, C2_30, X__dp[29], X__dn[29], Y__dp[29], Y__dn[29], C1_29, C2_29);
  SD2DigitCom_30 U24 (Z__dp[30], Z__dn[30], C2_30, C1_30);
endmodule

module SD2PureRBA_30_1 (Z__dp, Z__dn, X__dp, X__dn, Y__dp, Y__dn);
  output [31:1] Z__dp, Z__dn;
  input [30:1] X__dp, X__dn;
  input [30:1] Y__dp, Y__dn;
  wire C1_10;
  wire C1_11;
  wire C1_12;
  wire C1_13;
  wire C1_14;
  wire C1_15;
  wire C1_16;
  wire C1_17;
  wire C1_18;
  wire C1_19;
  wire C1_2;
  wire C1_20;
  wire C1_21;
  wire C1_22;
  wire C1_23;
  wire C1_24;
  wire C1_25;
  wire C1_26;
  wire C1_27;
  wire C1_28;
  wire C1_29;
  wire C1_3;
  wire C1_30;
  wire C1_31;
  wire C1_4;
  wire C1_5;
  wire C1_6;
  wire C1_7;
  wire C1_8;
  wire C1_9;
  wire C1i;
  wire C2_10;
  wire C2_11;
  wire C2_12;
  wire C2_13;
  wire C2_14;
  wire C2_15;
  wire C2_16;
  wire C2_17;
  wire C2_18;
  wire C2_19;
  wire C2_2;
  wire C2_20;
  wire C2_21;
  wire C2_22;
  wire C2_23;
  wire C2_24;
  wire C2_25;
  wire C2_26;
  wire C2_27;
  wire C2_28;
  wire C2_29;
  wire C2_3;
  wire C2_30;
  wire C2_31;
  wire C2_4;
  wire C2_5;
  wire C2_6;
  wire C2_7;
  wire C2_8;
  wire C2_9;
  wire C2i;
  UBZero_1_1 U0 (C1i);
  NUBZero_1_1 U1 (C2i);
  SD2DigitRBA_1 U2 (Z__dp[1], Z__dn[1], C1_2, C2_2, X__dp[1], X__dn[1], Y__dp[1], Y__dn[1], C1i, C2i);
  SD2DigitRBA_2 U3 (Z__dp[2], Z__dn[2], C1_3, C2_3, X__dp[2], X__dn[2], Y__dp[2], Y__dn[2], C1_2, C2_2);
  SD2DigitRBA_3 U4 (Z__dp[3], Z__dn[3], C1_4, C2_4, X__dp[3], X__dn[3], Y__dp[3], Y__dn[3], C1_3, C2_3);
  SD2DigitRBA_4 U5 (Z__dp[4], Z__dn[4], C1_5, C2_5, X__dp[4], X__dn[4], Y__dp[4], Y__dn[4], C1_4, C2_4);
  SD2DigitRBA_5 U6 (Z__dp[5], Z__dn[5], C1_6, C2_6, X__dp[5], X__dn[5], Y__dp[5], Y__dn[5], C1_5, C2_5);
  SD2DigitRBA_6 U7 (Z__dp[6], Z__dn[6], C1_7, C2_7, X__dp[6], X__dn[6], Y__dp[6], Y__dn[6], C1_6, C2_6);
  SD2DigitRBA_7 U8 (Z__dp[7], Z__dn[7], C1_8, C2_8, X__dp[7], X__dn[7], Y__dp[7], Y__dn[7], C1_7, C2_7);
  SD2DigitRBA_8 U9 (Z__dp[8], Z__dn[8], C1_9, C2_9, X__dp[8], X__dn[8], Y__dp[8], Y__dn[8], C1_8, C2_8);
  SD2DigitRBA_9 U10 (Z__dp[9], Z__dn[9], C1_10, C2_10, X__dp[9], X__dn[9], Y__dp[9], Y__dn[9], C1_9, C2_9);
  SD2DigitRBA_10 U11 (Z__dp[10], Z__dn[10], C1_11, C2_11, X__dp[10], X__dn[10], Y__dp[10], Y__dn[10], C1_10, C2_10);
  SD2DigitRBA_11 U12 (Z__dp[11], Z__dn[11], C1_12, C2_12, X__dp[11], X__dn[11], Y__dp[11], Y__dn[11], C1_11, C2_11);
  SD2DigitRBA_12 U13 (Z__dp[12], Z__dn[12], C1_13, C2_13, X__dp[12], X__dn[12], Y__dp[12], Y__dn[12], C1_12, C2_12);
  SD2DigitRBA_13 U14 (Z__dp[13], Z__dn[13], C1_14, C2_14, X__dp[13], X__dn[13], Y__dp[13], Y__dn[13], C1_13, C2_13);
  SD2DigitRBA_14 U15 (Z__dp[14], Z__dn[14], C1_15, C2_15, X__dp[14], X__dn[14], Y__dp[14], Y__dn[14], C1_14, C2_14);
  SD2DigitRBA_15 U16 (Z__dp[15], Z__dn[15], C1_16, C2_16, X__dp[15], X__dn[15], Y__dp[15], Y__dn[15], C1_15, C2_15);
  SD2DigitRBA_16 U17 (Z__dp[16], Z__dn[16], C1_17, C2_17, X__dp[16], X__dn[16], Y__dp[16], Y__dn[16], C1_16, C2_16);
  SD2DigitRBA_17 U18 (Z__dp[17], Z__dn[17], C1_18, C2_18, X__dp[17], X__dn[17], Y__dp[17], Y__dn[17], C1_17, C2_17);
  SD2DigitRBA_18 U19 (Z__dp[18], Z__dn[18], C1_19, C2_19, X__dp[18], X__dn[18], Y__dp[18], Y__dn[18], C1_18, C2_18);
  SD2DigitRBA_19 U20 (Z__dp[19], Z__dn[19], C1_20, C2_20, X__dp[19], X__dn[19], Y__dp[19], Y__dn[19], C1_19, C2_19);
  SD2DigitRBA_20 U21 (Z__dp[20], Z__dn[20], C1_21, C2_21, X__dp[20], X__dn[20], Y__dp[20], Y__dn[20], C1_20, C2_20);
  SD2DigitRBA_21 U22 (Z__dp[21], Z__dn[21], C1_22, C2_22, X__dp[21], X__dn[21], Y__dp[21], Y__dn[21], C1_21, C2_21);
  SD2DigitRBA_22 U23 (Z__dp[22], Z__dn[22], C1_23, C2_23, X__dp[22], X__dn[22], Y__dp[22], Y__dn[22], C1_22, C2_22);
  SD2DigitRBA_23 U24 (Z__dp[23], Z__dn[23], C1_24, C2_24, X__dp[23], X__dn[23], Y__dp[23], Y__dn[23], C1_23, C2_23);
  SD2DigitRBA_24 U25 (Z__dp[24], Z__dn[24], C1_25, C2_25, X__dp[24], X__dn[24], Y__dp[24], Y__dn[24], C1_24, C2_24);
  SD2DigitRBA_25 U26 (Z__dp[25], Z__dn[25], C1_26, C2_26, X__dp[25], X__dn[25], Y__dp[25], Y__dn[25], C1_25, C2_25);
  SD2DigitRBA_26 U27 (Z__dp[26], Z__dn[26], C1_27, C2_27, X__dp[26], X__dn[26], Y__dp[26], Y__dn[26], C1_26, C2_26);
  SD2DigitRBA_27 U28 (Z__dp[27], Z__dn[27], C1_28, C2_28, X__dp[27], X__dn[27], Y__dp[27], Y__dn[27], C1_27, C2_27);
  SD2DigitRBA_28 U29 (Z__dp[28], Z__dn[28], C1_29, C2_29, X__dp[28], X__dn[28], Y__dp[28], Y__dn[28], C1_28, C2_28);
  SD2DigitRBA_29 U30 (Z__dp[29], Z__dn[29], C1_30, C2_30, X__dp[29], X__dn[29], Y__dp[29], Y__dn[29], C1_29, C2_29);
  SD2DigitRBA_30 U31 (Z__dp[30], Z__dn[30], C1_31, C2_31, X__dp[30], X__dn[30], Y__dp[30], Y__dn[30], C1_30, C2_30);
  SD2DigitCom_31 U32 (Z__dp[31], Z__dn[31], C2_31, C1_31);
endmodule

module SD2RBA_16_0_18_2 (Z__dp, Z__dn, X__dp, X__dn, Y__dp, Y__dn);
  output [19:0] Z__dp, Z__dn;
  input [16:0] X__dp, X__dn;
  input [18:2] Y__dp, Y__dn;
  wire [18:0] XX__dp, XX__dn;
  wire [18:17] Zero__dp, Zero__dn;
  SD2_PN_A_Zero_18_000 U0 (Zero__dp[18:17], Zero__dn[18:17]);
  SD2_PN_ACMBIN_18_000 U1 (XX__dp[18:0], XX__dn[18:0], Zero__dp[18:17], Zero__dn[18:17], X__dp[16:0], X__dn[16:0]);
  SD2PureRBA_18_2 U2 (Z__dp[19:2], Z__dn[19:2], XX__dp[18:2], XX__dn[18:2], Y__dp[18:2], Y__dn[18:2]);
  SD2_PN_ACON_1_0 U3 (Z__dp[1:0], Z__dn[1:0], XX__dp[1:0], XX__dn[1:0]);
endmodule

module SD2RBA_19_0_23_4 (Z__dp, Z__dn, X__dp, X__dn, Y__dp, Y__dn);
  output [24:0] Z__dp, Z__dn;
  input [19:0] X__dp, X__dn;
  input [23:4] Y__dp, Y__dn;
  wire [23:0] XX__dp, XX__dn;
  wire [23:20] Zero__dp, Zero__dn;
  SD2_PN_A_Zero_23_000 U0 (Zero__dp[23:20], Zero__dn[23:20]);
  SD2_PN_ACMBIN_23_000 U1 (XX__dp[23:0], XX__dn[23:0], Zero__dp[23:20], Zero__dn[23:20], X__dp[19:0], X__dn[19:0]);
  SD2PureRBA_23_4 U2 (Z__dp[24:4], Z__dn[24:4], XX__dp[23:4], XX__dn[23:4], Y__dp[23:4], Y__dn[23:4]);
  SD2_PN_ACON_3_0 U3 (Z__dp[3:0], Z__dn[3:0], XX__dp[3:0], XX__dn[3:0]);
endmodule

module SD2RBA_20_4_22_6 (Z__dp, Z__dn, X__dp, X__dn, Y__dp, Y__dn);
  output [23:4] Z__dp, Z__dn;
  input [20:4] X__dp, X__dn;
  input [22:6] Y__dp, Y__dn;
  wire [22:4] XX__dp, XX__dn;
  wire [22:21] Zero__dp, Zero__dn;
  SD2_PN_A_Zero_22_000 U0 (Zero__dp[22:21], Zero__dn[22:21]);
  SD2_PN_ACMBIN_22_000 U1 (XX__dp[22:4], XX__dn[22:4], Zero__dp[22:21], Zero__dn[22:21], X__dp[20:4], X__dn[20:4]);
  SD2PureRBA_22_6 U2 (Z__dp[23:6], Z__dn[23:6], XX__dp[22:6], XX__dn[22:6], Y__dp[22:6], Y__dn[22:6]);
  SD2_PN_ACON_5_4 U3 (Z__dp[5:4], Z__dn[5:4], XX__dp[5:4], XX__dn[5:4]);
endmodule

module SD2RBA_24_0_30_1 (Z__dp, Z__dn, X__dp, X__dn, Y__dp, Y__dn);
  output [31:0] Z__dp, Z__dn;
  input [24:0] X__dp, X__dn;
  input [30:1] Y__dp, Y__dn;
  wire [30:0] XX__dp, XX__dn;
  wire [30:25] Zero__dp, Zero__dn;
  SD2_PN_A_Zero_30_000 U0 (Zero__dp[30:25], Zero__dn[30:25]);
  SD2_PN_ACMBIN_30_000 U1 (XX__dp[30:0], XX__dn[30:0], Zero__dp[30:25], Zero__dn[30:25], X__dp[24:0], X__dn[24:0]);
  SD2PureRBA_30_1 U2 (Z__dp[31:1], Z__dn[31:1], XX__dp[30:1], XX__dn[30:1], Y__dp[30:1], Y__dn[30:1]);
  SD2_PN_A1DCON_0 U3 (Z__dp[0], Z__dn[0], XX__dp[0], XX__dn[0]);
endmodule

module SD2RBA_24_8_26_10 (Z__dp, Z__dn, X__dp, X__dn, Y__dp, Y__dn);
  output [27:8] Z__dp, Z__dn;
  input [24:8] X__dp, X__dn;
  input [26:10] Y__dp, Y__dn;
  wire [26:8] XX__dp, XX__dn;
  wire [26:25] Zero__dp, Zero__dn;
  SD2_PN_A_Zero_26_000 U0 (Zero__dp[26:25], Zero__dn[26:25]);
  SD2_PN_ACMBIN_26_000 U1 (XX__dp[26:8], XX__dn[26:8], Zero__dp[26:25], Zero__dn[26:25], X__dp[24:8], X__dn[24:8]);
  SD2PureRBA_26_10 U2 (Z__dp[27:10], Z__dn[27:10], XX__dp[26:10], XX__dn[26:10], Y__dp[26:10], Y__dn[26:10]);
  SD2_PN_ACON_9_8 U3 (Z__dp[9:8], Z__dn[9:8], XX__dp[9:8], XX__dn[9:8]);
endmodule

module SD2RBA_27_8_29_1 (Z__dp, Z__dn, X__dp, X__dn, Y__dp, Y__dn);
  output [30:1] Z__dp, Z__dn;
  input [27:8] X__dp, X__dn;
  input [29:1] Y__dp, Y__dn;
  wire [29:8] XX__dp, XX__dn;
  wire [29:28] Zero__dp, Zero__dn;
  SD2_PN_A_Zero_29_000 U0 (Zero__dp[29:28], Zero__dn[29:28]);
  SD2_PN_ACMBIN_29_000 U1 (XX__dp[29:8], XX__dn[29:8], Zero__dp[29:28], Zero__dn[29:28], X__dp[27:8], X__dn[27:8]);
  SD2PureRBA_29_8 U2 (Z__dp[30:8], Z__dn[30:8], XX__dp[29:8], XX__dn[29:8], Y__dp[29:8], Y__dn[29:8]);
  SD2_PN_ACON_7_1 U3 (Z__dp[7:1], Z__dn[7:1], Y__dp[7:1], Y__dn[7:1]);
endmodule

module SD2RBA_28_12_28_1 (Z__dp, Z__dn, X__dp, X__dn, Y__dp, Y__dn);
  output [29:1] Z__dp, Z__dn;
  input [28:12] X__dp, X__dn;
  input [28:1] Y__dp, Y__dn;
  SD2PureRBA_28_12 U0 (Z__dp[29:12], Z__dn[29:12], X__dp[28:12], X__dn[28:12], Y__dp[28:12], Y__dn[28:12]);
  SD2_PN_ACON_11_1 U1 (Z__dp[11:1], Z__dn[11:1], Y__dp[11:1], Y__dn[11:1]);
endmodule

module SD2RBTR_16_0_18_2000 (Z__dp, Z__dn, PP0__dp, PP0__dn, PP1__dp, PP1__dn, PP2__dp, PP2__dn, PP3__dp, PP3__dn, PP4__dp, PP4__dn, PP5__dp, PP5__dn, PP6__dp, PP6__dn, PP7__dp, PP7__dn);
  output [31:0] Z__dp, Z__dn;
  input [16:0] PP0__dp, PP0__dn;
  input [18:2] PP1__dp, PP1__dn;
  input [20:4] PP2__dp, PP2__dn;
  input [22:6] PP3__dp, PP3__dn;
  input [24:8] PP4__dp, PP4__dn;
  input [26:10] PP5__dp, PP5__dn;
  input [28:12] PP6__dp, PP6__dn;
  input [28:1] PP7__dp, PP7__dn;
  wire [19:0] W1_0__dp, W1_0__dn;
  wire [23:4] W1_1__dp, W1_1__dn;
  wire [27:8] W1_2__dp, W1_2__dn;
  wire [29:1] W1_3__dp, W1_3__dn;
  wire [24:0] W2_4__dp, W2_4__dn;
  wire [30:1] W2_5__dp, W2_5__dn;
  SD2RBA_16_0_18_2 U0 (W1_0__dp[19:0], W1_0__dn[19:0], PP0__dp, PP0__dn, PP1__dp, PP1__dn);
  SD2RBA_20_4_22_6 U1 (W1_1__dp[23:4], W1_1__dn[23:4], PP2__dp, PP2__dn, PP3__dp, PP3__dn);
  SD2RBA_24_8_26_10 U2 (W1_2__dp[27:8], W1_2__dn[27:8], PP4__dp, PP4__dn, PP5__dp, PP5__dn);
  SD2RBA_28_12_28_1 U3 (W1_3__dp[29:1], W1_3__dn[29:1], PP6__dp, PP6__dn, PP7__dp, PP7__dn);
  SD2RBA_19_0_23_4 U4 (W2_4__dp[24:0], W2_4__dn[24:0], W1_0__dp[19:0], W1_0__dn[19:0], W1_1__dp[23:4], W1_1__dn[23:4]);
  SD2RBA_27_8_29_1 U5 (W2_5__dp[30:1], W2_5__dn[30:1], W1_2__dp[27:8], W1_2__dn[27:8], W1_3__dp[29:1], W1_3__dn[29:1]);
  SD2RBA_24_0_30_1 U6 (Z__dp[31:0], Z__dn[31:0], W2_4__dp[24:0], W2_4__dn[24:0], W2_5__dp[30:1], W2_5__dn[30:1]);
endmodule

module SD2TCConv_FCSkA_3000 (O, I__dp, I__dn);
  output [32:0] O;
  input [31:0] I__dp, I__dn;
  wire C;
  wire [32:0] S;
  wire [31:0] X;
  wire [31:0] Y;
  wire Z;
  SD2Decom_PN_31_0 U0 (X, Y, I__dp, I__dn);
  UBOne_0 U1 (C);
  UBPriFCSkA_31_0 U2 (S, X, Y, C);
  UBInv_32 U3 (Z, S[32]);
  TCCom_32_0 U4 (O, Z, S[31:0]);
endmodule

module SD2_PN_ACMBIN_18_000 (O__dp, O__dn, IN0__dp, IN0__dn, IN1__dp, IN1__dn);
  output [18:0] O__dp, O__dn;
  input [18:17] IN0__dp, IN0__dn;
  input [16:0] IN1__dp, IN1__dn;
  SD2_PN_ACON_18_17 U0 (O__dp[18:17], O__dn[18:17], IN0__dp, IN0__dn);
  SD2_PN_ACON_16_0 U1 (O__dp[16:0], O__dn[16:0], IN1__dp, IN1__dn);
endmodule

module SD2_PN_ACMBIN_22_000 (O__dp, O__dn, IN0__dp, IN0__dn, IN1__dp, IN1__dn);
  output [22:4] O__dp, O__dn;
  input [22:21] IN0__dp, IN0__dn;
  input [20:4] IN1__dp, IN1__dn;
  SD2_PN_ACON_22_21 U0 (O__dp[22:21], O__dn[22:21], IN0__dp, IN0__dn);
  SD2_PN_ACON_20_4 U1 (O__dp[20:4], O__dn[20:4], IN1__dp, IN1__dn);
endmodule

module SD2_PN_ACMBIN_23_000 (O__dp, O__dn, IN0__dp, IN0__dn, IN1__dp, IN1__dn);
  output [23:0] O__dp, O__dn;
  input [23:20] IN0__dp, IN0__dn;
  input [19:0] IN1__dp, IN1__dn;
  SD2_PN_ACON_23_20 U0 (O__dp[23:20], O__dn[23:20], IN0__dp, IN0__dn);
  SD2_PN_ACON_19_0 U1 (O__dp[19:0], O__dn[19:0], IN1__dp, IN1__dn);
endmodule

module SD2_PN_ACMBIN_26_000 (O__dp, O__dn, IN0__dp, IN0__dn, IN1__dp, IN1__dn);
  output [26:8] O__dp, O__dn;
  input [26:25] IN0__dp, IN0__dn;
  input [24:8] IN1__dp, IN1__dn;
  SD2_PN_ACON_26_25 U0 (O__dp[26:25], O__dn[26:25], IN0__dp, IN0__dn);
  SD2_PN_ACON_24_8 U1 (O__dp[24:8], O__dn[24:8], IN1__dp, IN1__dn);
endmodule

module SD2_PN_ACMBIN_29_000 (O__dp, O__dn, IN0__dp, IN0__dn, IN1__dp, IN1__dn);
  output [29:8] O__dp, O__dn;
  input [29:28] IN0__dp, IN0__dn;
  input [27:8] IN1__dp, IN1__dn;
  SD2_PN_ACON_29_28 U0 (O__dp[29:28], O__dn[29:28], IN0__dp, IN0__dn);
  SD2_PN_ACON_27_8 U1 (O__dp[27:8], O__dn[27:8], IN1__dp, IN1__dn);
endmodule

module SD2_PN_ACMBIN_30_000 (O__dp, O__dn, IN0__dp, IN0__dn, IN1__dp, IN1__dn);
  output [30:0] O__dp, O__dn;
  input [30:25] IN0__dp, IN0__dn;
  input [24:0] IN1__dp, IN1__dn;
  SD2_PN_ACON_30_25 U0 (O__dp[30:25], O__dn[30:25], IN0__dp, IN0__dn);
  SD2_PN_ACON_24_0 U1 (O__dp[24:0], O__dn[24:0], IN1__dp, IN1__dn);
endmodule

module SD2_PN_ACON_11_1 (O__dp, O__dn, I__dp, I__dn);
  output [11:1] O__dp, O__dn;
  input [11:1] I__dp, I__dn;
  SD2_PN_A1DCON_1 U0 (O__dp[1], O__dn[1], I__dp[1], I__dn[1]);
  SD2_PN_A1DCON_2 U1 (O__dp[2], O__dn[2], I__dp[2], I__dn[2]);
  SD2_PN_A1DCON_3 U2 (O__dp[3], O__dn[3], I__dp[3], I__dn[3]);
  SD2_PN_A1DCON_4 U3 (O__dp[4], O__dn[4], I__dp[4], I__dn[4]);
  SD2_PN_A1DCON_5 U4 (O__dp[5], O__dn[5], I__dp[5], I__dn[5]);
  SD2_PN_A1DCON_6 U5 (O__dp[6], O__dn[6], I__dp[6], I__dn[6]);
  SD2_PN_A1DCON_7 U6 (O__dp[7], O__dn[7], I__dp[7], I__dn[7]);
  SD2_PN_A1DCON_8 U7 (O__dp[8], O__dn[8], I__dp[8], I__dn[8]);
  SD2_PN_A1DCON_9 U8 (O__dp[9], O__dn[9], I__dp[9], I__dn[9]);
  SD2_PN_A1DCON_10 U9 (O__dp[10], O__dn[10], I__dp[10], I__dn[10]);
  SD2_PN_A1DCON_11 U10 (O__dp[11], O__dn[11], I__dp[11], I__dn[11]);
endmodule

module SD2_PN_ACON_16_0 (O__dp, O__dn, I__dp, I__dn);
  output [16:0] O__dp, O__dn;
  input [16:0] I__dp, I__dn;
  SD2_PN_A1DCON_0 U0 (O__dp[0], O__dn[0], I__dp[0], I__dn[0]);
  SD2_PN_A1DCON_1 U1 (O__dp[1], O__dn[1], I__dp[1], I__dn[1]);
  SD2_PN_A1DCON_2 U2 (O__dp[2], O__dn[2], I__dp[2], I__dn[2]);
  SD2_PN_A1DCON_3 U3 (O__dp[3], O__dn[3], I__dp[3], I__dn[3]);
  SD2_PN_A1DCON_4 U4 (O__dp[4], O__dn[4], I__dp[4], I__dn[4]);
  SD2_PN_A1DCON_5 U5 (O__dp[5], O__dn[5], I__dp[5], I__dn[5]);
  SD2_PN_A1DCON_6 U6 (O__dp[6], O__dn[6], I__dp[6], I__dn[6]);
  SD2_PN_A1DCON_7 U7 (O__dp[7], O__dn[7], I__dp[7], I__dn[7]);
  SD2_PN_A1DCON_8 U8 (O__dp[8], O__dn[8], I__dp[8], I__dn[8]);
  SD2_PN_A1DCON_9 U9 (O__dp[9], O__dn[9], I__dp[9], I__dn[9]);
  SD2_PN_A1DCON_10 U10 (O__dp[10], O__dn[10], I__dp[10], I__dn[10]);
  SD2_PN_A1DCON_11 U11 (O__dp[11], O__dn[11], I__dp[11], I__dn[11]);
  SD2_PN_A1DCON_12 U12 (O__dp[12], O__dn[12], I__dp[12], I__dn[12]);
  SD2_PN_A1DCON_13 U13 (O__dp[13], O__dn[13], I__dp[13], I__dn[13]);
  SD2_PN_A1DCON_14 U14 (O__dp[14], O__dn[14], I__dp[14], I__dn[14]);
  SD2_PN_A1DCON_15 U15 (O__dp[15], O__dn[15], I__dp[15], I__dn[15]);
  SD2_PN_A1DCON_16 U16 (O__dp[16], O__dn[16], I__dp[16], I__dn[16]);
endmodule

module SD2_PN_ACON_18_17 (O__dp, O__dn, I__dp, I__dn);
  output [18:17] O__dp, O__dn;
  input [18:17] I__dp, I__dn;
  SD2_PN_A1DCON_17 U0 (O__dp[17], O__dn[17], I__dp[17], I__dn[17]);
  SD2_PN_A1DCON_18 U1 (O__dp[18], O__dn[18], I__dp[18], I__dn[18]);
endmodule

module SD2_PN_ACON_19_0 (O__dp, O__dn, I__dp, I__dn);
  output [19:0] O__dp, O__dn;
  input [19:0] I__dp, I__dn;
  SD2_PN_A1DCON_0 U0 (O__dp[0], O__dn[0], I__dp[0], I__dn[0]);
  SD2_PN_A1DCON_1 U1 (O__dp[1], O__dn[1], I__dp[1], I__dn[1]);
  SD2_PN_A1DCON_2 U2 (O__dp[2], O__dn[2], I__dp[2], I__dn[2]);
  SD2_PN_A1DCON_3 U3 (O__dp[3], O__dn[3], I__dp[3], I__dn[3]);
  SD2_PN_A1DCON_4 U4 (O__dp[4], O__dn[4], I__dp[4], I__dn[4]);
  SD2_PN_A1DCON_5 U5 (O__dp[5], O__dn[5], I__dp[5], I__dn[5]);
  SD2_PN_A1DCON_6 U6 (O__dp[6], O__dn[6], I__dp[6], I__dn[6]);
  SD2_PN_A1DCON_7 U7 (O__dp[7], O__dn[7], I__dp[7], I__dn[7]);
  SD2_PN_A1DCON_8 U8 (O__dp[8], O__dn[8], I__dp[8], I__dn[8]);
  SD2_PN_A1DCON_9 U9 (O__dp[9], O__dn[9], I__dp[9], I__dn[9]);
  SD2_PN_A1DCON_10 U10 (O__dp[10], O__dn[10], I__dp[10], I__dn[10]);
  SD2_PN_A1DCON_11 U11 (O__dp[11], O__dn[11], I__dp[11], I__dn[11]);
  SD2_PN_A1DCON_12 U12 (O__dp[12], O__dn[12], I__dp[12], I__dn[12]);
  SD2_PN_A1DCON_13 U13 (O__dp[13], O__dn[13], I__dp[13], I__dn[13]);
  SD2_PN_A1DCON_14 U14 (O__dp[14], O__dn[14], I__dp[14], I__dn[14]);
  SD2_PN_A1DCON_15 U15 (O__dp[15], O__dn[15], I__dp[15], I__dn[15]);
  SD2_PN_A1DCON_16 U16 (O__dp[16], O__dn[16], I__dp[16], I__dn[16]);
  SD2_PN_A1DCON_17 U17 (O__dp[17], O__dn[17], I__dp[17], I__dn[17]);
  SD2_PN_A1DCON_18 U18 (O__dp[18], O__dn[18], I__dp[18], I__dn[18]);
  SD2_PN_A1DCON_19 U19 (O__dp[19], O__dn[19], I__dp[19], I__dn[19]);
endmodule

module SD2_PN_ACON_1_0 (O__dp, O__dn, I__dp, I__dn);
  output [1:0] O__dp, O__dn;
  input [1:0] I__dp, I__dn;
  SD2_PN_A1DCON_0 U0 (O__dp[0], O__dn[0], I__dp[0], I__dn[0]);
  SD2_PN_A1DCON_1 U1 (O__dp[1], O__dn[1], I__dp[1], I__dn[1]);
endmodule

module SD2_PN_ACON_20_4 (O__dp, O__dn, I__dp, I__dn);
  output [20:4] O__dp, O__dn;
  input [20:4] I__dp, I__dn;
  SD2_PN_A1DCON_4 U0 (O__dp[4], O__dn[4], I__dp[4], I__dn[4]);
  SD2_PN_A1DCON_5 U1 (O__dp[5], O__dn[5], I__dp[5], I__dn[5]);
  SD2_PN_A1DCON_6 U2 (O__dp[6], O__dn[6], I__dp[6], I__dn[6]);
  SD2_PN_A1DCON_7 U3 (O__dp[7], O__dn[7], I__dp[7], I__dn[7]);
  SD2_PN_A1DCON_8 U4 (O__dp[8], O__dn[8], I__dp[8], I__dn[8]);
  SD2_PN_A1DCON_9 U5 (O__dp[9], O__dn[9], I__dp[9], I__dn[9]);
  SD2_PN_A1DCON_10 U6 (O__dp[10], O__dn[10], I__dp[10], I__dn[10]);
  SD2_PN_A1DCON_11 U7 (O__dp[11], O__dn[11], I__dp[11], I__dn[11]);
  SD2_PN_A1DCON_12 U8 (O__dp[12], O__dn[12], I__dp[12], I__dn[12]);
  SD2_PN_A1DCON_13 U9 (O__dp[13], O__dn[13], I__dp[13], I__dn[13]);
  SD2_PN_A1DCON_14 U10 (O__dp[14], O__dn[14], I__dp[14], I__dn[14]);
  SD2_PN_A1DCON_15 U11 (O__dp[15], O__dn[15], I__dp[15], I__dn[15]);
  SD2_PN_A1DCON_16 U12 (O__dp[16], O__dn[16], I__dp[16], I__dn[16]);
  SD2_PN_A1DCON_17 U13 (O__dp[17], O__dn[17], I__dp[17], I__dn[17]);
  SD2_PN_A1DCON_18 U14 (O__dp[18], O__dn[18], I__dp[18], I__dn[18]);
  SD2_PN_A1DCON_19 U15 (O__dp[19], O__dn[19], I__dp[19], I__dn[19]);
  SD2_PN_A1DCON_20 U16 (O__dp[20], O__dn[20], I__dp[20], I__dn[20]);
endmodule

module SD2_PN_ACON_22_21 (O__dp, O__dn, I__dp, I__dn);
  output [22:21] O__dp, O__dn;
  input [22:21] I__dp, I__dn;
  SD2_PN_A1DCON_21 U0 (O__dp[21], O__dn[21], I__dp[21], I__dn[21]);
  SD2_PN_A1DCON_22 U1 (O__dp[22], O__dn[22], I__dp[22], I__dn[22]);
endmodule

module SD2_PN_ACON_23_20 (O__dp, O__dn, I__dp, I__dn);
  output [23:20] O__dp, O__dn;
  input [23:20] I__dp, I__dn;
  SD2_PN_A1DCON_20 U0 (O__dp[20], O__dn[20], I__dp[20], I__dn[20]);
  SD2_PN_A1DCON_21 U1 (O__dp[21], O__dn[21], I__dp[21], I__dn[21]);
  SD2_PN_A1DCON_22 U2 (O__dp[22], O__dn[22], I__dp[22], I__dn[22]);
  SD2_PN_A1DCON_23 U3 (O__dp[23], O__dn[23], I__dp[23], I__dn[23]);
endmodule

module SD2_PN_ACON_24_0 (O__dp, O__dn, I__dp, I__dn);
  output [24:0] O__dp, O__dn;
  input [24:0] I__dp, I__dn;
  SD2_PN_A1DCON_0 U0 (O__dp[0], O__dn[0], I__dp[0], I__dn[0]);
  SD2_PN_A1DCON_1 U1 (O__dp[1], O__dn[1], I__dp[1], I__dn[1]);
  SD2_PN_A1DCON_2 U2 (O__dp[2], O__dn[2], I__dp[2], I__dn[2]);
  SD2_PN_A1DCON_3 U3 (O__dp[3], O__dn[3], I__dp[3], I__dn[3]);
  SD2_PN_A1DCON_4 U4 (O__dp[4], O__dn[4], I__dp[4], I__dn[4]);
  SD2_PN_A1DCON_5 U5 (O__dp[5], O__dn[5], I__dp[5], I__dn[5]);
  SD2_PN_A1DCON_6 U6 (O__dp[6], O__dn[6], I__dp[6], I__dn[6]);
  SD2_PN_A1DCON_7 U7 (O__dp[7], O__dn[7], I__dp[7], I__dn[7]);
  SD2_PN_A1DCON_8 U8 (O__dp[8], O__dn[8], I__dp[8], I__dn[8]);
  SD2_PN_A1DCON_9 U9 (O__dp[9], O__dn[9], I__dp[9], I__dn[9]);
  SD2_PN_A1DCON_10 U10 (O__dp[10], O__dn[10], I__dp[10], I__dn[10]);
  SD2_PN_A1DCON_11 U11 (O__dp[11], O__dn[11], I__dp[11], I__dn[11]);
  SD2_PN_A1DCON_12 U12 (O__dp[12], O__dn[12], I__dp[12], I__dn[12]);
  SD2_PN_A1DCON_13 U13 (O__dp[13], O__dn[13], I__dp[13], I__dn[13]);
  SD2_PN_A1DCON_14 U14 (O__dp[14], O__dn[14], I__dp[14], I__dn[14]);
  SD2_PN_A1DCON_15 U15 (O__dp[15], O__dn[15], I__dp[15], I__dn[15]);
  SD2_PN_A1DCON_16 U16 (O__dp[16], O__dn[16], I__dp[16], I__dn[16]);
  SD2_PN_A1DCON_17 U17 (O__dp[17], O__dn[17], I__dp[17], I__dn[17]);
  SD2_PN_A1DCON_18 U18 (O__dp[18], O__dn[18], I__dp[18], I__dn[18]);
  SD2_PN_A1DCON_19 U19 (O__dp[19], O__dn[19], I__dp[19], I__dn[19]);
  SD2_PN_A1DCON_20 U20 (O__dp[20], O__dn[20], I__dp[20], I__dn[20]);
  SD2_PN_A1DCON_21 U21 (O__dp[21], O__dn[21], I__dp[21], I__dn[21]);
  SD2_PN_A1DCON_22 U22 (O__dp[22], O__dn[22], I__dp[22], I__dn[22]);
  SD2_PN_A1DCON_23 U23 (O__dp[23], O__dn[23], I__dp[23], I__dn[23]);
  SD2_PN_A1DCON_24 U24 (O__dp[24], O__dn[24], I__dp[24], I__dn[24]);
endmodule

module SD2_PN_ACON_24_8 (O__dp, O__dn, I__dp, I__dn);
  output [24:8] O__dp, O__dn;
  input [24:8] I__dp, I__dn;
  SD2_PN_A1DCON_8 U0 (O__dp[8], O__dn[8], I__dp[8], I__dn[8]);
  SD2_PN_A1DCON_9 U1 (O__dp[9], O__dn[9], I__dp[9], I__dn[9]);
  SD2_PN_A1DCON_10 U2 (O__dp[10], O__dn[10], I__dp[10], I__dn[10]);
  SD2_PN_A1DCON_11 U3 (O__dp[11], O__dn[11], I__dp[11], I__dn[11]);
  SD2_PN_A1DCON_12 U4 (O__dp[12], O__dn[12], I__dp[12], I__dn[12]);
  SD2_PN_A1DCON_13 U5 (O__dp[13], O__dn[13], I__dp[13], I__dn[13]);
  SD2_PN_A1DCON_14 U6 (O__dp[14], O__dn[14], I__dp[14], I__dn[14]);
  SD2_PN_A1DCON_15 U7 (O__dp[15], O__dn[15], I__dp[15], I__dn[15]);
  SD2_PN_A1DCON_16 U8 (O__dp[16], O__dn[16], I__dp[16], I__dn[16]);
  SD2_PN_A1DCON_17 U9 (O__dp[17], O__dn[17], I__dp[17], I__dn[17]);
  SD2_PN_A1DCON_18 U10 (O__dp[18], O__dn[18], I__dp[18], I__dn[18]);
  SD2_PN_A1DCON_19 U11 (O__dp[19], O__dn[19], I__dp[19], I__dn[19]);
  SD2_PN_A1DCON_20 U12 (O__dp[20], O__dn[20], I__dp[20], I__dn[20]);
  SD2_PN_A1DCON_21 U13 (O__dp[21], O__dn[21], I__dp[21], I__dn[21]);
  SD2_PN_A1DCON_22 U14 (O__dp[22], O__dn[22], I__dp[22], I__dn[22]);
  SD2_PN_A1DCON_23 U15 (O__dp[23], O__dn[23], I__dp[23], I__dn[23]);
  SD2_PN_A1DCON_24 U16 (O__dp[24], O__dn[24], I__dp[24], I__dn[24]);
endmodule

module SD2_PN_ACON_26_25 (O__dp, O__dn, I__dp, I__dn);
  output [26:25] O__dp, O__dn;
  input [26:25] I__dp, I__dn;
  SD2_PN_A1DCON_25 U0 (O__dp[25], O__dn[25], I__dp[25], I__dn[25]);
  SD2_PN_A1DCON_26 U1 (O__dp[26], O__dn[26], I__dp[26], I__dn[26]);
endmodule

module SD2_PN_ACON_27_8 (O__dp, O__dn, I__dp, I__dn);
  output [27:8] O__dp, O__dn;
  input [27:8] I__dp, I__dn;
  SD2_PN_A1DCON_8 U0 (O__dp[8], O__dn[8], I__dp[8], I__dn[8]);
  SD2_PN_A1DCON_9 U1 (O__dp[9], O__dn[9], I__dp[9], I__dn[9]);
  SD2_PN_A1DCON_10 U2 (O__dp[10], O__dn[10], I__dp[10], I__dn[10]);
  SD2_PN_A1DCON_11 U3 (O__dp[11], O__dn[11], I__dp[11], I__dn[11]);
  SD2_PN_A1DCON_12 U4 (O__dp[12], O__dn[12], I__dp[12], I__dn[12]);
  SD2_PN_A1DCON_13 U5 (O__dp[13], O__dn[13], I__dp[13], I__dn[13]);
  SD2_PN_A1DCON_14 U6 (O__dp[14], O__dn[14], I__dp[14], I__dn[14]);
  SD2_PN_A1DCON_15 U7 (O__dp[15], O__dn[15], I__dp[15], I__dn[15]);
  SD2_PN_A1DCON_16 U8 (O__dp[16], O__dn[16], I__dp[16], I__dn[16]);
  SD2_PN_A1DCON_17 U9 (O__dp[17], O__dn[17], I__dp[17], I__dn[17]);
  SD2_PN_A1DCON_18 U10 (O__dp[18], O__dn[18], I__dp[18], I__dn[18]);
  SD2_PN_A1DCON_19 U11 (O__dp[19], O__dn[19], I__dp[19], I__dn[19]);
  SD2_PN_A1DCON_20 U12 (O__dp[20], O__dn[20], I__dp[20], I__dn[20]);
  SD2_PN_A1DCON_21 U13 (O__dp[21], O__dn[21], I__dp[21], I__dn[21]);
  SD2_PN_A1DCON_22 U14 (O__dp[22], O__dn[22], I__dp[22], I__dn[22]);
  SD2_PN_A1DCON_23 U15 (O__dp[23], O__dn[23], I__dp[23], I__dn[23]);
  SD2_PN_A1DCON_24 U16 (O__dp[24], O__dn[24], I__dp[24], I__dn[24]);
  SD2_PN_A1DCON_25 U17 (O__dp[25], O__dn[25], I__dp[25], I__dn[25]);
  SD2_PN_A1DCON_26 U18 (O__dp[26], O__dn[26], I__dp[26], I__dn[26]);
  SD2_PN_A1DCON_27 U19 (O__dp[27], O__dn[27], I__dp[27], I__dn[27]);
endmodule

module SD2_PN_ACON_29_28 (O__dp, O__dn, I__dp, I__dn);
  output [29:28] O__dp, O__dn;
  input [29:28] I__dp, I__dn;
  SD2_PN_A1DCON_28 U0 (O__dp[28], O__dn[28], I__dp[28], I__dn[28]);
  SD2_PN_A1DCON_29 U1 (O__dp[29], O__dn[29], I__dp[29], I__dn[29]);
endmodule

module SD2_PN_ACON_30_25 (O__dp, O__dn, I__dp, I__dn);
  output [30:25] O__dp, O__dn;
  input [30:25] I__dp, I__dn;
  SD2_PN_A1DCON_25 U0 (O__dp[25], O__dn[25], I__dp[25], I__dn[25]);
  SD2_PN_A1DCON_26 U1 (O__dp[26], O__dn[26], I__dp[26], I__dn[26]);
  SD2_PN_A1DCON_27 U2 (O__dp[27], O__dn[27], I__dp[27], I__dn[27]);
  SD2_PN_A1DCON_28 U3 (O__dp[28], O__dn[28], I__dp[28], I__dn[28]);
  SD2_PN_A1DCON_29 U4 (O__dp[29], O__dn[29], I__dp[29], I__dn[29]);
  SD2_PN_A1DCON_30 U5 (O__dp[30], O__dn[30], I__dp[30], I__dn[30]);
endmodule

module SD2_PN_ACON_3_0 (O__dp, O__dn, I__dp, I__dn);
  output [3:0] O__dp, O__dn;
  input [3:0] I__dp, I__dn;
  SD2_PN_A1DCON_0 U0 (O__dp[0], O__dn[0], I__dp[0], I__dn[0]);
  SD2_PN_A1DCON_1 U1 (O__dp[1], O__dn[1], I__dp[1], I__dn[1]);
  SD2_PN_A1DCON_2 U2 (O__dp[2], O__dn[2], I__dp[2], I__dn[2]);
  SD2_PN_A1DCON_3 U3 (O__dp[3], O__dn[3], I__dp[3], I__dn[3]);
endmodule

module SD2_PN_ACON_5_4 (O__dp, O__dn, I__dp, I__dn);
  output [5:4] O__dp, O__dn;
  input [5:4] I__dp, I__dn;
  SD2_PN_A1DCON_4 U0 (O__dp[4], O__dn[4], I__dp[4], I__dn[4]);
  SD2_PN_A1DCON_5 U1 (O__dp[5], O__dn[5], I__dp[5], I__dn[5]);
endmodule

module SD2_PN_ACON_7_1 (O__dp, O__dn, I__dp, I__dn);
  output [7:1] O__dp, O__dn;
  input [7:1] I__dp, I__dn;
  SD2_PN_A1DCON_1 U0 (O__dp[1], O__dn[1], I__dp[1], I__dn[1]);
  SD2_PN_A1DCON_2 U1 (O__dp[2], O__dn[2], I__dp[2], I__dn[2]);
  SD2_PN_A1DCON_3 U2 (O__dp[3], O__dn[3], I__dp[3], I__dn[3]);
  SD2_PN_A1DCON_4 U3 (O__dp[4], O__dn[4], I__dp[4], I__dn[4]);
  SD2_PN_A1DCON_5 U4 (O__dp[5], O__dn[5], I__dp[5], I__dn[5]);
  SD2_PN_A1DCON_6 U5 (O__dp[6], O__dn[6], I__dp[6], I__dn[6]);
  SD2_PN_A1DCON_7 U6 (O__dp[7], O__dn[7], I__dp[7], I__dn[7]);
endmodule

module SD2_PN_ACON_9_8 (O__dp, O__dn, I__dp, I__dn);
  output [9:8] O__dp, O__dn;
  input [9:8] I__dp, I__dn;
  SD2_PN_A1DCON_8 U0 (O__dp[8], O__dn[8], I__dp[8], I__dn[8]);
  SD2_PN_A1DCON_9 U1 (O__dp[9], O__dn[9], I__dp[9], I__dn[9]);
endmodule

module UBCMBIN_16_16_14_000 (O, IN0, IN1);
  output [16:0] O;
  input IN0;
  input [14:0] IN1;
  UB1DCON_16 U0 (O[16], IN0);
  UBZero_15_15 U1 (O[15]);
  UBCON_14_0 U2 (O[14:0], IN1);
endmodule

module UBCMBIN_18_18_16_000 (O, IN0, IN1);
  output [18:2] O;
  input IN0;
  input [16:2] IN1;
  UB1DCON_18 U0 (O[18], IN0);
  UBZero_17_17 U1 (O[17]);
  UBCON_16_2 U2 (O[16:2], IN1);
endmodule

module UBCMBIN_20_20_18_000 (O, IN0, IN1);
  output [20:4] O;
  input IN0;
  input [18:4] IN1;
  UB1DCON_20 U0 (O[20], IN0);
  UBZero_19_19 U1 (O[19]);
  UBCON_18_4 U2 (O[18:4], IN1);
endmodule

module UBCMBIN_22_22_20_000 (O, IN0, IN1);
  output [22:6] O;
  input IN0;
  input [20:6] IN1;
  UB1DCON_22 U0 (O[22], IN0);
  UBZero_21_21 U1 (O[21]);
  UBCON_20_6 U2 (O[20:6], IN1);
endmodule

module UBCMBIN_24_24_22_000 (O, IN0, IN1);
  output [24:8] O;
  input IN0;
  input [22:8] IN1;
  UB1DCON_24 U0 (O[24], IN0);
  UBZero_23_23 U1 (O[23]);
  UBCON_22_8 U2 (O[22:8], IN1);
endmodule

module UBCMBIN_26_26_24_000 (O, IN0, IN1);
  output [26:10] O;
  input IN0;
  input [24:10] IN1;
  UB1DCON_26 U0 (O[26], IN0);
  UBZero_25_25 U1 (O[25]);
  UBCON_24_10 U2 (O[24:10], IN1);
endmodule

module UBCMBIN_28_14_13_000 (O, IN0, IN1);
  output [28:1] O;
  input [28:14] IN0;
  input [13:1] IN1;
  UBCON_28_14 U0 (O[28:14], IN0);
  UBCON_13_1 U1 (O[13:1], IN1);
endmodule

module UBCMBIN_28_28_26_000 (O, IN0, IN1);
  output [28:12] O;
  input IN0;
  input [26:12] IN1;
  UB1DCON_28 U0 (O[28], IN0);
  UBZero_27_27 U1 (O[27]);
  UBCON_26_12 U2 (O[26:12], IN1);
endmodule

module UBCON_13_1 (O, I);
  output [13:1] O;
  input [13:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
  UB1DCON_6 U5 (O[6], I[6]);
  UB1DCON_7 U6 (O[7], I[7]);
  UB1DCON_8 U7 (O[8], I[8]);
  UB1DCON_9 U8 (O[9], I[9]);
  UB1DCON_10 U9 (O[10], I[10]);
  UB1DCON_11 U10 (O[11], I[11]);
  UB1DCON_12 U11 (O[12], I[12]);
  UB1DCON_13 U12 (O[13], I[13]);
endmodule

module UBCON_14_0 (O, I);
  output [14:0] O;
  input [14:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
  UB1DCON_13 U13 (O[13], I[13]);
  UB1DCON_14 U14 (O[14], I[14]);
endmodule

module UBCON_16_2 (O, I);
  output [16:2] O;
  input [16:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
  UB1DCON_6 U4 (O[6], I[6]);
  UB1DCON_7 U5 (O[7], I[7]);
  UB1DCON_8 U6 (O[8], I[8]);
  UB1DCON_9 U7 (O[9], I[9]);
  UB1DCON_10 U8 (O[10], I[10]);
  UB1DCON_11 U9 (O[11], I[11]);
  UB1DCON_12 U10 (O[12], I[12]);
  UB1DCON_13 U11 (O[13], I[13]);
  UB1DCON_14 U12 (O[14], I[14]);
  UB1DCON_15 U13 (O[15], I[15]);
  UB1DCON_16 U14 (O[16], I[16]);
endmodule

module UBCON_18_4 (O, I);
  output [18:4] O;
  input [18:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
  UB1DCON_11 U7 (O[11], I[11]);
  UB1DCON_12 U8 (O[12], I[12]);
  UB1DCON_13 U9 (O[13], I[13]);
  UB1DCON_14 U10 (O[14], I[14]);
  UB1DCON_15 U11 (O[15], I[15]);
  UB1DCON_16 U12 (O[16], I[16]);
  UB1DCON_17 U13 (O[17], I[17]);
  UB1DCON_18 U14 (O[18], I[18]);
endmodule

module UBCON_20_6 (O, I);
  output [20:6] O;
  input [20:6] I;
  UB1DCON_6 U0 (O[6], I[6]);
  UB1DCON_7 U1 (O[7], I[7]);
  UB1DCON_8 U2 (O[8], I[8]);
  UB1DCON_9 U3 (O[9], I[9]);
  UB1DCON_10 U4 (O[10], I[10]);
  UB1DCON_11 U5 (O[11], I[11]);
  UB1DCON_12 U6 (O[12], I[12]);
  UB1DCON_13 U7 (O[13], I[13]);
  UB1DCON_14 U8 (O[14], I[14]);
  UB1DCON_15 U9 (O[15], I[15]);
  UB1DCON_16 U10 (O[16], I[16]);
  UB1DCON_17 U11 (O[17], I[17]);
  UB1DCON_18 U12 (O[18], I[18]);
  UB1DCON_19 U13 (O[19], I[19]);
  UB1DCON_20 U14 (O[20], I[20]);
endmodule

module UBCON_22_8 (O, I);
  output [22:8] O;
  input [22:8] I;
  UB1DCON_8 U0 (O[8], I[8]);
  UB1DCON_9 U1 (O[9], I[9]);
  UB1DCON_10 U2 (O[10], I[10]);
  UB1DCON_11 U3 (O[11], I[11]);
  UB1DCON_12 U4 (O[12], I[12]);
  UB1DCON_13 U5 (O[13], I[13]);
  UB1DCON_14 U6 (O[14], I[14]);
  UB1DCON_15 U7 (O[15], I[15]);
  UB1DCON_16 U8 (O[16], I[16]);
  UB1DCON_17 U9 (O[17], I[17]);
  UB1DCON_18 U10 (O[18], I[18]);
  UB1DCON_19 U11 (O[19], I[19]);
  UB1DCON_20 U12 (O[20], I[20]);
  UB1DCON_21 U13 (O[21], I[21]);
  UB1DCON_22 U14 (O[22], I[22]);
endmodule

module UBCON_24_10 (O, I);
  output [24:10] O;
  input [24:10] I;
  UB1DCON_10 U0 (O[10], I[10]);
  UB1DCON_11 U1 (O[11], I[11]);
  UB1DCON_12 U2 (O[12], I[12]);
  UB1DCON_13 U3 (O[13], I[13]);
  UB1DCON_14 U4 (O[14], I[14]);
  UB1DCON_15 U5 (O[15], I[15]);
  UB1DCON_16 U6 (O[16], I[16]);
  UB1DCON_17 U7 (O[17], I[17]);
  UB1DCON_18 U8 (O[18], I[18]);
  UB1DCON_19 U9 (O[19], I[19]);
  UB1DCON_20 U10 (O[20], I[20]);
  UB1DCON_21 U11 (O[21], I[21]);
  UB1DCON_22 U12 (O[22], I[22]);
  UB1DCON_23 U13 (O[23], I[23]);
  UB1DCON_24 U14 (O[24], I[24]);
endmodule

module UBCON_26_12 (O, I);
  output [26:12] O;
  input [26:12] I;
  UB1DCON_12 U0 (O[12], I[12]);
  UB1DCON_13 U1 (O[13], I[13]);
  UB1DCON_14 U2 (O[14], I[14]);
  UB1DCON_15 U3 (O[15], I[15]);
  UB1DCON_16 U4 (O[16], I[16]);
  UB1DCON_17 U5 (O[17], I[17]);
  UB1DCON_18 U6 (O[18], I[18]);
  UB1DCON_19 U7 (O[19], I[19]);
  UB1DCON_20 U8 (O[20], I[20]);
  UB1DCON_21 U9 (O[21], I[21]);
  UB1DCON_22 U10 (O[22], I[22]);
  UB1DCON_23 U11 (O[23], I[23]);
  UB1DCON_24 U12 (O[24], I[24]);
  UB1DCON_25 U13 (O[25], I[25]);
  UB1DCON_26 U14 (O[26], I[26]);
endmodule

module UBCON_28_14 (O, I);
  output [28:14] O;
  input [28:14] I;
  UB1DCON_14 U0 (O[14], I[14]);
  UB1DCON_15 U1 (O[15], I[15]);
  UB1DCON_16 U2 (O[16], I[16]);
  UB1DCON_17 U3 (O[17], I[17]);
  UB1DCON_18 U4 (O[18], I[18]);
  UB1DCON_19 U5 (O[19], I[19]);
  UB1DCON_20 U6 (O[20], I[20]);
  UB1DCON_21 U7 (O[21], I[21]);
  UB1DCON_22 U8 (O[22], I[22]);
  UB1DCON_23 U9 (O[23], I[23]);
  UB1DCON_24 U10 (O[24], I[24]);
  UB1DCON_25 U11 (O[25], I[25]);
  UB1DCON_26 U12 (O[26], I[26]);
  UB1DCON_27 U13 (O[27], I[27]);
  UB1DCON_28 U14 (O[28], I[28]);
endmodule

module UBMinusVPPG_14_0_000 (P, PP, C, I1, I2);
  output C;
  output P;
  output [15:1] PP;
  input [14:0] I1;
  input I2;
  wire S;
  wire [15:1] W;
  UB1BPPG_0_1 U0 (W[1], I1[0], I2);
  UB1BPPG_1_1 U1 (W[2], I1[1], I2);
  UB1BPPG_2_1 U2 (W[3], I1[2], I2);
  UB1BPPG_3_1 U3 (W[4], I1[3], I2);
  UB1BPPG_4_1 U4 (W[5], I1[4], I2);
  UB1BPPG_5_1 U5 (W[6], I1[5], I2);
  UB1BPPG_6_1 U6 (W[7], I1[6], I2);
  UB1BPPG_7_1 U7 (W[8], I1[7], I2);
  UB1BPPG_8_1 U8 (W[9], I1[8], I2);
  UB1BPPG_9_1 U9 (W[10], I1[9], I2);
  UB1BPPG_10_1 U10 (W[11], I1[10], I2);
  UB1BPPG_11_1 U11 (W[12], I1[11], I2);
  UB1BPPG_12_1 U12 (W[13], I1[12], I2);
  UB1BPPG_13_1 U13 (W[14], I1[13], I2);
  UB1BPPG_14_1 U14 (W[15], I1[14], I2);
  SignP_0 U15 (S);
  UBNUBWCON_15_1 U16 (PP, W, S);
  NUBBBG_1 U17 (C, S);
  UBHBBG_16 U18 (P, S);
endmodule

module UBMinusVPPG_14_0_001 (P, PP, C, I1, I2);
  output C;
  output P;
  output [17:3] PP;
  input [14:0] I1;
  input I2;
  wire S;
  wire [17:3] W;
  UB1BPPG_0_3 U0 (W[3], I1[0], I2);
  UB1BPPG_1_3 U1 (W[4], I1[1], I2);
  UB1BPPG_2_3 U2 (W[5], I1[2], I2);
  UB1BPPG_3_3 U3 (W[6], I1[3], I2);
  UB1BPPG_4_3 U4 (W[7], I1[4], I2);
  UB1BPPG_5_3 U5 (W[8], I1[5], I2);
  UB1BPPG_6_3 U6 (W[9], I1[6], I2);
  UB1BPPG_7_3 U7 (W[10], I1[7], I2);
  UB1BPPG_8_3 U8 (W[11], I1[8], I2);
  UB1BPPG_9_3 U9 (W[12], I1[9], I2);
  UB1BPPG_10_3 U10 (W[13], I1[10], I2);
  UB1BPPG_11_3 U11 (W[14], I1[11], I2);
  UB1BPPG_12_3 U12 (W[15], I1[12], I2);
  UB1BPPG_13_3 U13 (W[16], I1[13], I2);
  UB1BPPG_14_3 U14 (W[17], I1[14], I2);
  SignP_0 U15 (S);
  UBNUBWCON_17_3 U16 (PP, W, S);
  NUBBBG_3 U17 (C, S);
  UBHBBG_18 U18 (P, S);
endmodule

module UBMinusVPPG_14_0_002 (P, PP, C, I1, I2);
  output C;
  output P;
  output [19:5] PP;
  input [14:0] I1;
  input I2;
  wire S;
  wire [19:5] W;
  UB1BPPG_0_5 U0 (W[5], I1[0], I2);
  UB1BPPG_1_5 U1 (W[6], I1[1], I2);
  UB1BPPG_2_5 U2 (W[7], I1[2], I2);
  UB1BPPG_3_5 U3 (W[8], I1[3], I2);
  UB1BPPG_4_5 U4 (W[9], I1[4], I2);
  UB1BPPG_5_5 U5 (W[10], I1[5], I2);
  UB1BPPG_6_5 U6 (W[11], I1[6], I2);
  UB1BPPG_7_5 U7 (W[12], I1[7], I2);
  UB1BPPG_8_5 U8 (W[13], I1[8], I2);
  UB1BPPG_9_5 U9 (W[14], I1[9], I2);
  UB1BPPG_10_5 U10 (W[15], I1[10], I2);
  UB1BPPG_11_5 U11 (W[16], I1[11], I2);
  UB1BPPG_12_5 U12 (W[17], I1[12], I2);
  UB1BPPG_13_5 U13 (W[18], I1[13], I2);
  UB1BPPG_14_5 U14 (W[19], I1[14], I2);
  SignP_0 U15 (S);
  UBNUBWCON_19_5 U16 (PP, W, S);
  NUBBBG_5 U17 (C, S);
  UBHBBG_20 U18 (P, S);
endmodule

module UBMinusVPPG_14_0_003 (P, PP, C, I1, I2);
  output C;
  output P;
  output [21:7] PP;
  input [14:0] I1;
  input I2;
  wire S;
  wire [21:7] W;
  UB1BPPG_0_7 U0 (W[7], I1[0], I2);
  UB1BPPG_1_7 U1 (W[8], I1[1], I2);
  UB1BPPG_2_7 U2 (W[9], I1[2], I2);
  UB1BPPG_3_7 U3 (W[10], I1[3], I2);
  UB1BPPG_4_7 U4 (W[11], I1[4], I2);
  UB1BPPG_5_7 U5 (W[12], I1[5], I2);
  UB1BPPG_6_7 U6 (W[13], I1[6], I2);
  UB1BPPG_7_7 U7 (W[14], I1[7], I2);
  UB1BPPG_8_7 U8 (W[15], I1[8], I2);
  UB1BPPG_9_7 U9 (W[16], I1[9], I2);
  UB1BPPG_10_7 U10 (W[17], I1[10], I2);
  UB1BPPG_11_7 U11 (W[18], I1[11], I2);
  UB1BPPG_12_7 U12 (W[19], I1[12], I2);
  UB1BPPG_13_7 U13 (W[20], I1[13], I2);
  UB1BPPG_14_7 U14 (W[21], I1[14], I2);
  SignP_0 U15 (S);
  UBNUBWCON_21_7 U16 (PP, W, S);
  NUBBBG_7 U17 (C, S);
  UBHBBG_22 U18 (P, S);
endmodule

module UBMinusVPPG_14_0_004 (P, PP, C, I1, I2);
  output C;
  output P;
  output [23:9] PP;
  input [14:0] I1;
  input I2;
  wire S;
  wire [23:9] W;
  UB1BPPG_0_9 U0 (W[9], I1[0], I2);
  UB1BPPG_1_9 U1 (W[10], I1[1], I2);
  UB1BPPG_2_9 U2 (W[11], I1[2], I2);
  UB1BPPG_3_9 U3 (W[12], I1[3], I2);
  UB1BPPG_4_9 U4 (W[13], I1[4], I2);
  UB1BPPG_5_9 U5 (W[14], I1[5], I2);
  UB1BPPG_6_9 U6 (W[15], I1[6], I2);
  UB1BPPG_7_9 U7 (W[16], I1[7], I2);
  UB1BPPG_8_9 U8 (W[17], I1[8], I2);
  UB1BPPG_9_9 U9 (W[18], I1[9], I2);
  UB1BPPG_10_9 U10 (W[19], I1[10], I2);
  UB1BPPG_11_9 U11 (W[20], I1[11], I2);
  UB1BPPG_12_9 U12 (W[21], I1[12], I2);
  UB1BPPG_13_9 U13 (W[22], I1[13], I2);
  UB1BPPG_14_9 U14 (W[23], I1[14], I2);
  SignP_0 U15 (S);
  UBNUBWCON_23_9 U16 (PP, W, S);
  NUBBBG_9 U17 (C, S);
  UBHBBG_24 U18 (P, S);
endmodule

module UBMinusVPPG_14_0_005 (P, PP, C, I1, I2);
  output C;
  output P;
  output [25:11] PP;
  input [14:0] I1;
  input I2;
  wire S;
  wire [25:11] W;
  UB1BPPG_0_11 U0 (W[11], I1[0], I2);
  UB1BPPG_1_11 U1 (W[12], I1[1], I2);
  UB1BPPG_2_11 U2 (W[13], I1[2], I2);
  UB1BPPG_3_11 U3 (W[14], I1[3], I2);
  UB1BPPG_4_11 U4 (W[15], I1[4], I2);
  UB1BPPG_5_11 U5 (W[16], I1[5], I2);
  UB1BPPG_6_11 U6 (W[17], I1[6], I2);
  UB1BPPG_7_11 U7 (W[18], I1[7], I2);
  UB1BPPG_8_11 U8 (W[19], I1[8], I2);
  UB1BPPG_9_11 U9 (W[20], I1[9], I2);
  UB1BPPG_10_11 U10 (W[21], I1[10], I2);
  UB1BPPG_11_11 U11 (W[22], I1[11], I2);
  UB1BPPG_12_11 U12 (W[23], I1[12], I2);
  UB1BPPG_13_11 U13 (W[24], I1[13], I2);
  UB1BPPG_14_11 U14 (W[25], I1[14], I2);
  SignP_0 U15 (S);
  UBNUBWCON_25_11 U16 (PP, W, S);
  NUBBBG_11 U17 (C, S);
  UBHBBG_26 U18 (P, S);
endmodule

module UBMinusVPPG_14_0_006 (P, PP, C, I1, I2);
  output C;
  output P;
  output [27:13] PP;
  input [14:0] I1;
  input I2;
  wire S;
  wire [27:13] W;
  UB1BPPG_0_13 U0 (W[13], I1[0], I2);
  UB1BPPG_1_13 U1 (W[14], I1[1], I2);
  UB1BPPG_2_13 U2 (W[15], I1[2], I2);
  UB1BPPG_3_13 U3 (W[16], I1[3], I2);
  UB1BPPG_4_13 U4 (W[17], I1[4], I2);
  UB1BPPG_5_13 U5 (W[18], I1[5], I2);
  UB1BPPG_6_13 U6 (W[19], I1[6], I2);
  UB1BPPG_7_13 U7 (W[20], I1[7], I2);
  UB1BPPG_8_13 U8 (W[21], I1[8], I2);
  UB1BPPG_9_13 U9 (W[22], I1[9], I2);
  UB1BPPG_10_13 U10 (W[23], I1[10], I2);
  UB1BPPG_11_13 U11 (W[24], I1[11], I2);
  UB1BPPG_12_13 U12 (W[25], I1[12], I2);
  UB1BPPG_13_13 U13 (W[26], I1[13], I2);
  UB1BPPG_14_13 U14 (W[27], I1[14], I2);
  SignP_0 U15 (S);
  UBNUBWCON_27_13 U16 (PP, W, S);
  NUBBBG_13 U17 (C, S);
  UBHBBG_28 U18 (P, S);
endmodule

module UBNUBWCON_15_1 (O, I, S);
  output [15:1] O;
  input [15:1] I;
  input S;
  BWCPN_1 U0 (O[1], I[1], S);
  BWCPN_2 U1 (O[2], I[2], S);
  BWCPN_3 U2 (O[3], I[3], S);
  BWCPN_4 U3 (O[4], I[4], S);
  BWCPN_5 U4 (O[5], I[5], S);
  BWCPN_6 U5 (O[6], I[6], S);
  BWCPN_7 U6 (O[7], I[7], S);
  BWCPN_8 U7 (O[8], I[8], S);
  BWCPN_9 U8 (O[9], I[9], S);
  BWCPN_10 U9 (O[10], I[10], S);
  BWCPN_11 U10 (O[11], I[11], S);
  BWCPN_12 U11 (O[12], I[12], S);
  BWCPN_13 U12 (O[13], I[13], S);
  BWCPN_14 U13 (O[14], I[14], S);
  BWCPN_15 U14 (O[15], I[15], S);
endmodule

module UBNUBWCON_17_3 (O, I, S);
  output [17:3] O;
  input [17:3] I;
  input S;
  BWCPN_3 U0 (O[3], I[3], S);
  BWCPN_4 U1 (O[4], I[4], S);
  BWCPN_5 U2 (O[5], I[5], S);
  BWCPN_6 U3 (O[6], I[6], S);
  BWCPN_7 U4 (O[7], I[7], S);
  BWCPN_8 U5 (O[8], I[8], S);
  BWCPN_9 U6 (O[9], I[9], S);
  BWCPN_10 U7 (O[10], I[10], S);
  BWCPN_11 U8 (O[11], I[11], S);
  BWCPN_12 U9 (O[12], I[12], S);
  BWCPN_13 U10 (O[13], I[13], S);
  BWCPN_14 U11 (O[14], I[14], S);
  BWCPN_15 U12 (O[15], I[15], S);
  BWCPN_16 U13 (O[16], I[16], S);
  BWCPN_17 U14 (O[17], I[17], S);
endmodule

module UBNUBWCON_19_5 (O, I, S);
  output [19:5] O;
  input [19:5] I;
  input S;
  BWCPN_5 U0 (O[5], I[5], S);
  BWCPN_6 U1 (O[6], I[6], S);
  BWCPN_7 U2 (O[7], I[7], S);
  BWCPN_8 U3 (O[8], I[8], S);
  BWCPN_9 U4 (O[9], I[9], S);
  BWCPN_10 U5 (O[10], I[10], S);
  BWCPN_11 U6 (O[11], I[11], S);
  BWCPN_12 U7 (O[12], I[12], S);
  BWCPN_13 U8 (O[13], I[13], S);
  BWCPN_14 U9 (O[14], I[14], S);
  BWCPN_15 U10 (O[15], I[15], S);
  BWCPN_16 U11 (O[16], I[16], S);
  BWCPN_17 U12 (O[17], I[17], S);
  BWCPN_18 U13 (O[18], I[18], S);
  BWCPN_19 U14 (O[19], I[19], S);
endmodule

module UBNUBWCON_21_7 (O, I, S);
  output [21:7] O;
  input [21:7] I;
  input S;
  BWCPN_7 U0 (O[7], I[7], S);
  BWCPN_8 U1 (O[8], I[8], S);
  BWCPN_9 U2 (O[9], I[9], S);
  BWCPN_10 U3 (O[10], I[10], S);
  BWCPN_11 U4 (O[11], I[11], S);
  BWCPN_12 U5 (O[12], I[12], S);
  BWCPN_13 U6 (O[13], I[13], S);
  BWCPN_14 U7 (O[14], I[14], S);
  BWCPN_15 U8 (O[15], I[15], S);
  BWCPN_16 U9 (O[16], I[16], S);
  BWCPN_17 U10 (O[17], I[17], S);
  BWCPN_18 U11 (O[18], I[18], S);
  BWCPN_19 U12 (O[19], I[19], S);
  BWCPN_20 U13 (O[20], I[20], S);
  BWCPN_21 U14 (O[21], I[21], S);
endmodule

module UBNUBWCON_23_9 (O, I, S);
  output [23:9] O;
  input [23:9] I;
  input S;
  BWCPN_9 U0 (O[9], I[9], S);
  BWCPN_10 U1 (O[10], I[10], S);
  BWCPN_11 U2 (O[11], I[11], S);
  BWCPN_12 U3 (O[12], I[12], S);
  BWCPN_13 U4 (O[13], I[13], S);
  BWCPN_14 U5 (O[14], I[14], S);
  BWCPN_15 U6 (O[15], I[15], S);
  BWCPN_16 U7 (O[16], I[16], S);
  BWCPN_17 U8 (O[17], I[17], S);
  BWCPN_18 U9 (O[18], I[18], S);
  BWCPN_19 U10 (O[19], I[19], S);
  BWCPN_20 U11 (O[20], I[20], S);
  BWCPN_21 U12 (O[21], I[21], S);
  BWCPN_22 U13 (O[22], I[22], S);
  BWCPN_23 U14 (O[23], I[23], S);
endmodule

module UBNUBWCON_25_11 (O, I, S);
  output [25:11] O;
  input [25:11] I;
  input S;
  BWCPN_11 U0 (O[11], I[11], S);
  BWCPN_12 U1 (O[12], I[12], S);
  BWCPN_13 U2 (O[13], I[13], S);
  BWCPN_14 U3 (O[14], I[14], S);
  BWCPN_15 U4 (O[15], I[15], S);
  BWCPN_16 U5 (O[16], I[16], S);
  BWCPN_17 U6 (O[17], I[17], S);
  BWCPN_18 U7 (O[18], I[18], S);
  BWCPN_19 U8 (O[19], I[19], S);
  BWCPN_20 U9 (O[20], I[20], S);
  BWCPN_21 U10 (O[21], I[21], S);
  BWCPN_22 U11 (O[22], I[22], S);
  BWCPN_23 U12 (O[23], I[23], S);
  BWCPN_24 U13 (O[24], I[24], S);
  BWCPN_25 U14 (O[25], I[25], S);
endmodule

module UBNUBWCON_27_13 (O, I, S);
  output [27:13] O;
  input [27:13] I;
  input S;
  BWCPN_13 U0 (O[13], I[13], S);
  BWCPN_14 U1 (O[14], I[14], S);
  BWCPN_15 U2 (O[15], I[15], S);
  BWCPN_16 U3 (O[16], I[16], S);
  BWCPN_17 U4 (O[17], I[17], S);
  BWCPN_18 U5 (O[18], I[18], S);
  BWCPN_19 U6 (O[19], I[19], S);
  BWCPN_20 U7 (O[20], I[20], S);
  BWCPN_21 U8 (O[21], I[21], S);
  BWCPN_22 U9 (O[22], I[22], S);
  BWCPN_23 U10 (O[23], I[23], S);
  BWCPN_24 U11 (O[24], I[24], S);
  BWCPN_25 U12 (O[25], I[25], S);
  BWCPN_26 U13 (O[26], I[26], S);
  BWCPN_27 U14 (O[27], I[27], S);
endmodule

module UBNUB_SD2Comp_16_000 (O__dp, O__dn, I_p, I_n);
  output [16:0] O__dp, O__dn;
  input [15:1] I_n;
  input [16:0] I_p;
  wire [16:0] N;
  wire Z_h;
  wire Z_l;
  NUBZero_16_16 U0 (Z_h);
  NUBZero_0_0 U1 (Z_l);
  NUBCMBIN_16_16_15000 U2 (N, Z_h, I_n, Z_l);
  UBNUB_SD2PriComp_000 U3 (O__dp, O__dn, I_p, N);
endmodule

module UBNUB_SD2Comp_18_000 (O__dp, O__dn, I_p, I_n);
  output [18:2] O__dp, O__dn;
  input [17:3] I_n;
  input [18:2] I_p;
  wire [18:2] N;
  wire Z_h;
  wire Z_l;
  NUBZero_18_18 U0 (Z_h);
  NUBZero_2_2 U1 (Z_l);
  NUBCMBIN_18_18_17000 U2 (N, Z_h, I_n, Z_l);
  UBNUB_SD2PriComp_001 U3 (O__dp, O__dn, I_p, N);
endmodule

module UBNUB_SD2Comp_20_000 (O__dp, O__dn, I_p, I_n);
  output [20:4] O__dp, O__dn;
  input [19:5] I_n;
  input [20:4] I_p;
  wire [20:4] N;
  wire Z_h;
  wire Z_l;
  NUBZero_20_20 U0 (Z_h);
  NUBZero_4_4 U1 (Z_l);
  NUBCMBIN_20_20_19000 U2 (N, Z_h, I_n, Z_l);
  UBNUB_SD2PriComp_002 U3 (O__dp, O__dn, I_p, N);
endmodule

module UBNUB_SD2Comp_22_000 (O__dp, O__dn, I_p, I_n);
  output [22:6] O__dp, O__dn;
  input [21:7] I_n;
  input [22:6] I_p;
  wire [22:6] N;
  wire Z_h;
  wire Z_l;
  NUBZero_22_22 U0 (Z_h);
  NUBZero_6_6 U1 (Z_l);
  NUBCMBIN_22_22_21000 U2 (N, Z_h, I_n, Z_l);
  UBNUB_SD2PriComp_003 U3 (O__dp, O__dn, I_p, N);
endmodule

module UBNUB_SD2Comp_24_000 (O__dp, O__dn, I_p, I_n);
  output [24:8] O__dp, O__dn;
  input [23:9] I_n;
  input [24:8] I_p;
  wire [24:8] N;
  wire Z_h;
  wire Z_l;
  NUBZero_24_24 U0 (Z_h);
  NUBZero_8_8 U1 (Z_l);
  NUBCMBIN_24_24_23000 U2 (N, Z_h, I_n, Z_l);
  UBNUB_SD2PriComp_004 U3 (O__dp, O__dn, I_p, N);
endmodule

module UBNUB_SD2Comp_26_000 (O__dp, O__dn, I_p, I_n);
  output [26:10] O__dp, O__dn;
  input [25:11] I_n;
  input [26:10] I_p;
  wire [26:10] N;
  wire Z_h;
  wire Z_l;
  NUBZero_26_26 U0 (Z_h);
  NUBZero_10_10 U1 (Z_l);
  NUBCMBIN_26_26_25000 U2 (N, Z_h, I_n, Z_l);
  UBNUB_SD2PriComp_005 U3 (O__dp, O__dn, I_p, N);
endmodule

module UBNUB_SD2Comp_28_000 (O__dp, O__dn, I_p, I_n);
  output [28:12] O__dp, O__dn;
  input [27:13] I_n;
  input [28:12] I_p;
  wire [28:12] N;
  wire Z_h;
  wire Z_l;
  NUBZero_28_28 U0 (Z_h);
  NUBZero_12_12 U1 (Z_l);
  NUBCMBIN_28_28_27000 U2 (N, Z_h, I_n, Z_l);
  UBNUB_SD2PriComp_006 U3 (O__dp, O__dn, I_p, N);
endmodule

module UBNUB_SD2Comp_28_001 (O__dp, O__dn, I_p, I_n);
  output [28:1] O__dp, O__dn;
  input [13:1] I_n;
  input [28:14] I_p;
  wire [28:1] N;
  wire [28:1] P;
  wire [28:14] Z_h;
  wire [13:1] Z_l;
  NUBZero_28_14 U0 (Z_h);
  UBZero_13_1 U1 (Z_l);
  UBCMBIN_28_14_13_000 U2 (P, I_p, Z_l);
  NUBCMBIN_28_14_13000 U3 (N, Z_h, I_n);
  UBNUB_SD2PriComp_007 U4 (O__dp, O__dn, P, N);
endmodule

module UBNUB_SD2PriComp_000 (O__dp, O__dn, I_p, I_n);
  output [16:0] O__dp, O__dn;
  input [16:0] I_n;
  input [16:0] I_p;
  SD2DigitCom_0 U0 (O__dp[0], O__dn[0], I_n[0], I_p[0]);
  SD2DigitCom_1 U1 (O__dp[1], O__dn[1], I_n[1], I_p[1]);
  SD2DigitCom_2 U2 (O__dp[2], O__dn[2], I_n[2], I_p[2]);
  SD2DigitCom_3 U3 (O__dp[3], O__dn[3], I_n[3], I_p[3]);
  SD2DigitCom_4 U4 (O__dp[4], O__dn[4], I_n[4], I_p[4]);
  SD2DigitCom_5 U5 (O__dp[5], O__dn[5], I_n[5], I_p[5]);
  SD2DigitCom_6 U6 (O__dp[6], O__dn[6], I_n[6], I_p[6]);
  SD2DigitCom_7 U7 (O__dp[7], O__dn[7], I_n[7], I_p[7]);
  SD2DigitCom_8 U8 (O__dp[8], O__dn[8], I_n[8], I_p[8]);
  SD2DigitCom_9 U9 (O__dp[9], O__dn[9], I_n[9], I_p[9]);
  SD2DigitCom_10 U10 (O__dp[10], O__dn[10], I_n[10], I_p[10]);
  SD2DigitCom_11 U11 (O__dp[11], O__dn[11], I_n[11], I_p[11]);
  SD2DigitCom_12 U12 (O__dp[12], O__dn[12], I_n[12], I_p[12]);
  SD2DigitCom_13 U13 (O__dp[13], O__dn[13], I_n[13], I_p[13]);
  SD2DigitCom_14 U14 (O__dp[14], O__dn[14], I_n[14], I_p[14]);
  SD2DigitCom_15 U15 (O__dp[15], O__dn[15], I_n[15], I_p[15]);
  SD2DigitCom_16 U16 (O__dp[16], O__dn[16], I_n[16], I_p[16]);
endmodule

module UBNUB_SD2PriComp_001 (O__dp, O__dn, I_p, I_n);
  output [18:2] O__dp, O__dn;
  input [18:2] I_n;
  input [18:2] I_p;
  SD2DigitCom_2 U0 (O__dp[2], O__dn[2], I_n[2], I_p[2]);
  SD2DigitCom_3 U1 (O__dp[3], O__dn[3], I_n[3], I_p[3]);
  SD2DigitCom_4 U2 (O__dp[4], O__dn[4], I_n[4], I_p[4]);
  SD2DigitCom_5 U3 (O__dp[5], O__dn[5], I_n[5], I_p[5]);
  SD2DigitCom_6 U4 (O__dp[6], O__dn[6], I_n[6], I_p[6]);
  SD2DigitCom_7 U5 (O__dp[7], O__dn[7], I_n[7], I_p[7]);
  SD2DigitCom_8 U6 (O__dp[8], O__dn[8], I_n[8], I_p[8]);
  SD2DigitCom_9 U7 (O__dp[9], O__dn[9], I_n[9], I_p[9]);
  SD2DigitCom_10 U8 (O__dp[10], O__dn[10], I_n[10], I_p[10]);
  SD2DigitCom_11 U9 (O__dp[11], O__dn[11], I_n[11], I_p[11]);
  SD2DigitCom_12 U10 (O__dp[12], O__dn[12], I_n[12], I_p[12]);
  SD2DigitCom_13 U11 (O__dp[13], O__dn[13], I_n[13], I_p[13]);
  SD2DigitCom_14 U12 (O__dp[14], O__dn[14], I_n[14], I_p[14]);
  SD2DigitCom_15 U13 (O__dp[15], O__dn[15], I_n[15], I_p[15]);
  SD2DigitCom_16 U14 (O__dp[16], O__dn[16], I_n[16], I_p[16]);
  SD2DigitCom_17 U15 (O__dp[17], O__dn[17], I_n[17], I_p[17]);
  SD2DigitCom_18 U16 (O__dp[18], O__dn[18], I_n[18], I_p[18]);
endmodule

module UBNUB_SD2PriComp_002 (O__dp, O__dn, I_p, I_n);
  output [20:4] O__dp, O__dn;
  input [20:4] I_n;
  input [20:4] I_p;
  SD2DigitCom_4 U0 (O__dp[4], O__dn[4], I_n[4], I_p[4]);
  SD2DigitCom_5 U1 (O__dp[5], O__dn[5], I_n[5], I_p[5]);
  SD2DigitCom_6 U2 (O__dp[6], O__dn[6], I_n[6], I_p[6]);
  SD2DigitCom_7 U3 (O__dp[7], O__dn[7], I_n[7], I_p[7]);
  SD2DigitCom_8 U4 (O__dp[8], O__dn[8], I_n[8], I_p[8]);
  SD2DigitCom_9 U5 (O__dp[9], O__dn[9], I_n[9], I_p[9]);
  SD2DigitCom_10 U6 (O__dp[10], O__dn[10], I_n[10], I_p[10]);
  SD2DigitCom_11 U7 (O__dp[11], O__dn[11], I_n[11], I_p[11]);
  SD2DigitCom_12 U8 (O__dp[12], O__dn[12], I_n[12], I_p[12]);
  SD2DigitCom_13 U9 (O__dp[13], O__dn[13], I_n[13], I_p[13]);
  SD2DigitCom_14 U10 (O__dp[14], O__dn[14], I_n[14], I_p[14]);
  SD2DigitCom_15 U11 (O__dp[15], O__dn[15], I_n[15], I_p[15]);
  SD2DigitCom_16 U12 (O__dp[16], O__dn[16], I_n[16], I_p[16]);
  SD2DigitCom_17 U13 (O__dp[17], O__dn[17], I_n[17], I_p[17]);
  SD2DigitCom_18 U14 (O__dp[18], O__dn[18], I_n[18], I_p[18]);
  SD2DigitCom_19 U15 (O__dp[19], O__dn[19], I_n[19], I_p[19]);
  SD2DigitCom_20 U16 (O__dp[20], O__dn[20], I_n[20], I_p[20]);
endmodule

module UBNUB_SD2PriComp_003 (O__dp, O__dn, I_p, I_n);
  output [22:6] O__dp, O__dn;
  input [22:6] I_n;
  input [22:6] I_p;
  SD2DigitCom_6 U0 (O__dp[6], O__dn[6], I_n[6], I_p[6]);
  SD2DigitCom_7 U1 (O__dp[7], O__dn[7], I_n[7], I_p[7]);
  SD2DigitCom_8 U2 (O__dp[8], O__dn[8], I_n[8], I_p[8]);
  SD2DigitCom_9 U3 (O__dp[9], O__dn[9], I_n[9], I_p[9]);
  SD2DigitCom_10 U4 (O__dp[10], O__dn[10], I_n[10], I_p[10]);
  SD2DigitCom_11 U5 (O__dp[11], O__dn[11], I_n[11], I_p[11]);
  SD2DigitCom_12 U6 (O__dp[12], O__dn[12], I_n[12], I_p[12]);
  SD2DigitCom_13 U7 (O__dp[13], O__dn[13], I_n[13], I_p[13]);
  SD2DigitCom_14 U8 (O__dp[14], O__dn[14], I_n[14], I_p[14]);
  SD2DigitCom_15 U9 (O__dp[15], O__dn[15], I_n[15], I_p[15]);
  SD2DigitCom_16 U10 (O__dp[16], O__dn[16], I_n[16], I_p[16]);
  SD2DigitCom_17 U11 (O__dp[17], O__dn[17], I_n[17], I_p[17]);
  SD2DigitCom_18 U12 (O__dp[18], O__dn[18], I_n[18], I_p[18]);
  SD2DigitCom_19 U13 (O__dp[19], O__dn[19], I_n[19], I_p[19]);
  SD2DigitCom_20 U14 (O__dp[20], O__dn[20], I_n[20], I_p[20]);
  SD2DigitCom_21 U15 (O__dp[21], O__dn[21], I_n[21], I_p[21]);
  SD2DigitCom_22 U16 (O__dp[22], O__dn[22], I_n[22], I_p[22]);
endmodule

module UBNUB_SD2PriComp_004 (O__dp, O__dn, I_p, I_n);
  output [24:8] O__dp, O__dn;
  input [24:8] I_n;
  input [24:8] I_p;
  SD2DigitCom_8 U0 (O__dp[8], O__dn[8], I_n[8], I_p[8]);
  SD2DigitCom_9 U1 (O__dp[9], O__dn[9], I_n[9], I_p[9]);
  SD2DigitCom_10 U2 (O__dp[10], O__dn[10], I_n[10], I_p[10]);
  SD2DigitCom_11 U3 (O__dp[11], O__dn[11], I_n[11], I_p[11]);
  SD2DigitCom_12 U4 (O__dp[12], O__dn[12], I_n[12], I_p[12]);
  SD2DigitCom_13 U5 (O__dp[13], O__dn[13], I_n[13], I_p[13]);
  SD2DigitCom_14 U6 (O__dp[14], O__dn[14], I_n[14], I_p[14]);
  SD2DigitCom_15 U7 (O__dp[15], O__dn[15], I_n[15], I_p[15]);
  SD2DigitCom_16 U8 (O__dp[16], O__dn[16], I_n[16], I_p[16]);
  SD2DigitCom_17 U9 (O__dp[17], O__dn[17], I_n[17], I_p[17]);
  SD2DigitCom_18 U10 (O__dp[18], O__dn[18], I_n[18], I_p[18]);
  SD2DigitCom_19 U11 (O__dp[19], O__dn[19], I_n[19], I_p[19]);
  SD2DigitCom_20 U12 (O__dp[20], O__dn[20], I_n[20], I_p[20]);
  SD2DigitCom_21 U13 (O__dp[21], O__dn[21], I_n[21], I_p[21]);
  SD2DigitCom_22 U14 (O__dp[22], O__dn[22], I_n[22], I_p[22]);
  SD2DigitCom_23 U15 (O__dp[23], O__dn[23], I_n[23], I_p[23]);
  SD2DigitCom_24 U16 (O__dp[24], O__dn[24], I_n[24], I_p[24]);
endmodule

module UBNUB_SD2PriComp_005 (O__dp, O__dn, I_p, I_n);
  output [26:10] O__dp, O__dn;
  input [26:10] I_n;
  input [26:10] I_p;
  SD2DigitCom_10 U0 (O__dp[10], O__dn[10], I_n[10], I_p[10]);
  SD2DigitCom_11 U1 (O__dp[11], O__dn[11], I_n[11], I_p[11]);
  SD2DigitCom_12 U2 (O__dp[12], O__dn[12], I_n[12], I_p[12]);
  SD2DigitCom_13 U3 (O__dp[13], O__dn[13], I_n[13], I_p[13]);
  SD2DigitCom_14 U4 (O__dp[14], O__dn[14], I_n[14], I_p[14]);
  SD2DigitCom_15 U5 (O__dp[15], O__dn[15], I_n[15], I_p[15]);
  SD2DigitCom_16 U6 (O__dp[16], O__dn[16], I_n[16], I_p[16]);
  SD2DigitCom_17 U7 (O__dp[17], O__dn[17], I_n[17], I_p[17]);
  SD2DigitCom_18 U8 (O__dp[18], O__dn[18], I_n[18], I_p[18]);
  SD2DigitCom_19 U9 (O__dp[19], O__dn[19], I_n[19], I_p[19]);
  SD2DigitCom_20 U10 (O__dp[20], O__dn[20], I_n[20], I_p[20]);
  SD2DigitCom_21 U11 (O__dp[21], O__dn[21], I_n[21], I_p[21]);
  SD2DigitCom_22 U12 (O__dp[22], O__dn[22], I_n[22], I_p[22]);
  SD2DigitCom_23 U13 (O__dp[23], O__dn[23], I_n[23], I_p[23]);
  SD2DigitCom_24 U14 (O__dp[24], O__dn[24], I_n[24], I_p[24]);
  SD2DigitCom_25 U15 (O__dp[25], O__dn[25], I_n[25], I_p[25]);
  SD2DigitCom_26 U16 (O__dp[26], O__dn[26], I_n[26], I_p[26]);
endmodule

module UBNUB_SD2PriComp_006 (O__dp, O__dn, I_p, I_n);
  output [28:12] O__dp, O__dn;
  input [28:12] I_n;
  input [28:12] I_p;
  SD2DigitCom_12 U0 (O__dp[12], O__dn[12], I_n[12], I_p[12]);
  SD2DigitCom_13 U1 (O__dp[13], O__dn[13], I_n[13], I_p[13]);
  SD2DigitCom_14 U2 (O__dp[14], O__dn[14], I_n[14], I_p[14]);
  SD2DigitCom_15 U3 (O__dp[15], O__dn[15], I_n[15], I_p[15]);
  SD2DigitCom_16 U4 (O__dp[16], O__dn[16], I_n[16], I_p[16]);
  SD2DigitCom_17 U5 (O__dp[17], O__dn[17], I_n[17], I_p[17]);
  SD2DigitCom_18 U6 (O__dp[18], O__dn[18], I_n[18], I_p[18]);
  SD2DigitCom_19 U7 (O__dp[19], O__dn[19], I_n[19], I_p[19]);
  SD2DigitCom_20 U8 (O__dp[20], O__dn[20], I_n[20], I_p[20]);
  SD2DigitCom_21 U9 (O__dp[21], O__dn[21], I_n[21], I_p[21]);
  SD2DigitCom_22 U10 (O__dp[22], O__dn[22], I_n[22], I_p[22]);
  SD2DigitCom_23 U11 (O__dp[23], O__dn[23], I_n[23], I_p[23]);
  SD2DigitCom_24 U12 (O__dp[24], O__dn[24], I_n[24], I_p[24]);
  SD2DigitCom_25 U13 (O__dp[25], O__dn[25], I_n[25], I_p[25]);
  SD2DigitCom_26 U14 (O__dp[26], O__dn[26], I_n[26], I_p[26]);
  SD2DigitCom_27 U15 (O__dp[27], O__dn[27], I_n[27], I_p[27]);
  SD2DigitCom_28 U16 (O__dp[28], O__dn[28], I_n[28], I_p[28]);
endmodule

module UBNUB_SD2PriComp_007 (O__dp, O__dn, I_p, I_n);
  output [28:1] O__dp, O__dn;
  input [28:1] I_n;
  input [28:1] I_p;
  SD2DigitCom_1 U0 (O__dp[1], O__dn[1], I_n[1], I_p[1]);
  SD2DigitCom_2 U1 (O__dp[2], O__dn[2], I_n[2], I_p[2]);
  SD2DigitCom_3 U2 (O__dp[3], O__dn[3], I_n[3], I_p[3]);
  SD2DigitCom_4 U3 (O__dp[4], O__dn[4], I_n[4], I_p[4]);
  SD2DigitCom_5 U4 (O__dp[5], O__dn[5], I_n[5], I_p[5]);
  SD2DigitCom_6 U5 (O__dp[6], O__dn[6], I_n[6], I_p[6]);
  SD2DigitCom_7 U6 (O__dp[7], O__dn[7], I_n[7], I_p[7]);
  SD2DigitCom_8 U7 (O__dp[8], O__dn[8], I_n[8], I_p[8]);
  SD2DigitCom_9 U8 (O__dp[9], O__dn[9], I_n[9], I_p[9]);
  SD2DigitCom_10 U9 (O__dp[10], O__dn[10], I_n[10], I_p[10]);
  SD2DigitCom_11 U10 (O__dp[11], O__dn[11], I_n[11], I_p[11]);
  SD2DigitCom_12 U11 (O__dp[12], O__dn[12], I_n[12], I_p[12]);
  SD2DigitCom_13 U12 (O__dp[13], O__dn[13], I_n[13], I_p[13]);
  SD2DigitCom_14 U13 (O__dp[14], O__dn[14], I_n[14], I_p[14]);
  SD2DigitCom_15 U14 (O__dp[15], O__dn[15], I_n[15], I_p[15]);
  SD2DigitCom_16 U15 (O__dp[16], O__dn[16], I_n[16], I_p[16]);
  SD2DigitCom_17 U16 (O__dp[17], O__dn[17], I_n[17], I_p[17]);
  SD2DigitCom_18 U17 (O__dp[18], O__dn[18], I_n[18], I_p[18]);
  SD2DigitCom_19 U18 (O__dp[19], O__dn[19], I_n[19], I_p[19]);
  SD2DigitCom_20 U19 (O__dp[20], O__dn[20], I_n[20], I_p[20]);
  SD2DigitCom_21 U20 (O__dp[21], O__dn[21], I_n[21], I_p[21]);
  SD2DigitCom_22 U21 (O__dp[22], O__dn[22], I_n[22], I_p[22]);
  SD2DigitCom_23 U22 (O__dp[23], O__dn[23], I_n[23], I_p[23]);
  SD2DigitCom_24 U23 (O__dp[24], O__dn[24], I_n[24], I_p[24]);
  SD2DigitCom_25 U24 (O__dp[25], O__dn[25], I_n[25], I_p[25]);
  SD2DigitCom_26 U25 (O__dp[26], O__dn[26], I_n[26], I_p[26]);
  SD2DigitCom_27 U26 (O__dp[27], O__dn[27], I_n[27], I_p[27]);
  SD2DigitCom_28 U27 (O__dp[28], O__dn[28], I_n[28], I_p[28]);
endmodule

module UBSPPG_14_0_14_0 (PP0__dp, PP0__dn, PP1__dp, PP1__dn, PP2__dp, PP2__dn, PP3__dp, PP3__dn, PP4__dp, PP4__dn, PP5__dp, PP5__dn, PP6__dp, PP6__dn, PP7__dp, PP7__dn, I1, I2);
  output [16:0] PP0__dp, PP0__dn;
  output [18:2] PP1__dp, PP1__dn;
  output [20:4] PP2__dp, PP2__dn;
  output [22:6] PP3__dp, PP3__dn;
  output [24:8] PP4__dp, PP4__dn;
  output [26:10] PP5__dp, PP5__dn;
  output [28:12] PP6__dp, PP6__dn;
  output [28:1] PP7__dp, PP7__dn;
  input [14:0] I1;
  input [14:0] I2;
  wire [13:1] MI_B;
  wire NCO0;
  wire NCO1;
  wire NCO2;
  wire NCO3;
  wire NCO4;
  wire NCO5;
  wire NCO6;
  wire [15:1] NPP0;
  wire [17:3] NPP1;
  wire [19:5] NPP2;
  wire [21:7] NPP3;
  wire [23:9] NPP4;
  wire [25:11] NPP5;
  wire [27:13] NPP6;
  wire POG0;
  wire POG1;
  wire POG2;
  wire POG3;
  wire POG4;
  wire POG5;
  wire POG6;
  wire [14:0] PPP0;
  wire [16:2] PPP1;
  wire [18:4] PPP2;
  wire [20:6] PPP3;
  wire [22:8] PPP4;
  wire [24:10] PPP5;
  wire [26:12] PPP6;
  wire [28:14] PPP7;
  wire [16:0] PP_p0;
  wire [18:2] PP_p1;
  wire [20:4] PP_p2;
  wire [22:6] PP_p3;
  wire [24:8] PP_p4;
  wire [26:10] PP_p5;
  wire [28:12] PP_p6;
  UBVPPG_14_0_0 U0 (PPP0, I1, I2[0]);
  UBMinusVPPG_14_0_000 U1 (POG0, NPP0, NCO0, I1, I2[1]);
  UBCMBIN_16_16_14_000 U2 (PP_p0, POG0, PPP0);
  UBNUB_SD2Comp_16_000 U3 (PP0__dp[16:0], PP0__dn[16:0], PP_p0, NPP0);
  UBVPPG_14_0_2 U4 (PPP1, I1, I2[2]);
  UBMinusVPPG_14_0_001 U5 (POG1, NPP1, NCO1, I1, I2[3]);
  UBCMBIN_18_18_16_000 U6 (PP_p1, POG1, PPP1);
  UBNUB_SD2Comp_18_000 U7 (PP1__dp[18:2], PP1__dn[18:2], PP_p1, NPP1);
  UBVPPG_14_0_4 U8 (PPP2, I1, I2[4]);
  UBMinusVPPG_14_0_002 U9 (POG2, NPP2, NCO2, I1, I2[5]);
  UBCMBIN_20_20_18_000 U10 (PP_p2, POG2, PPP2);
  UBNUB_SD2Comp_20_000 U11 (PP2__dp[20:4], PP2__dn[20:4], PP_p2, NPP2);
  UBVPPG_14_0_6 U12 (PPP3, I1, I2[6]);
  UBMinusVPPG_14_0_003 U13 (POG3, NPP3, NCO3, I1, I2[7]);
  UBCMBIN_22_22_20_000 U14 (PP_p3, POG3, PPP3);
  UBNUB_SD2Comp_22_000 U15 (PP3__dp[22:6], PP3__dn[22:6], PP_p3, NPP3);
  UBVPPG_14_0_8 U16 (PPP4, I1, I2[8]);
  UBMinusVPPG_14_0_004 U17 (POG4, NPP4, NCO4, I1, I2[9]);
  UBCMBIN_24_24_22_000 U18 (PP_p4, POG4, PPP4);
  UBNUB_SD2Comp_24_000 U19 (PP4__dp[24:8], PP4__dn[24:8], PP_p4, NPP4);
  UBVPPG_14_0_10 U20 (PPP5, I1, I2[10]);
  UBMinusVPPG_14_0_005 U21 (POG5, NPP5, NCO5, I1, I2[11]);
  UBCMBIN_26_26_24_000 U22 (PP_p5, POG5, PPP5);
  UBNUB_SD2Comp_26_000 U23 (PP5__dp[26:10], PP5__dn[26:10], PP_p5, NPP5);
  UBVPPG_14_0_12 U24 (PPP6, I1, I2[12]);
  UBMinusVPPG_14_0_006 U25 (POG6, NPP6, NCO6, I1, I2[13]);
  UBCMBIN_28_28_26_000 U26 (PP_p6, POG6, PPP6);
  UBNUB_SD2Comp_28_000 U27 (PP6__dp[28:12], PP6__dn[28:12], PP_p6, NPP6);
  NUBCMBIN_13_13_11000 U28 (MI_B, NCO6, NCO5, NCO4, NCO3, NCO2, NCO1, NCO0);
  UBVPPG_14_0_14 U29 (PPP7, I1, I2[14]);
  UBNUB_SD2Comp_28_001 U30 (PP7__dp[28:1], PP7__dn[28:1], PPP7, MI_B);
endmodule

module UBVPPG_14_0_0 (O, IN1, IN2);
  output [14:0] O;
  input [14:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
  UB1BPPG_6_0 U6 (O[6], IN1[6], IN2);
  UB1BPPG_7_0 U7 (O[7], IN1[7], IN2);
  UB1BPPG_8_0 U8 (O[8], IN1[8], IN2);
  UB1BPPG_9_0 U9 (O[9], IN1[9], IN2);
  UB1BPPG_10_0 U10 (O[10], IN1[10], IN2);
  UB1BPPG_11_0 U11 (O[11], IN1[11], IN2);
  UB1BPPG_12_0 U12 (O[12], IN1[12], IN2);
  UB1BPPG_13_0 U13 (O[13], IN1[13], IN2);
  UB1BPPG_14_0 U14 (O[14], IN1[14], IN2);
endmodule

module UBVPPG_14_0_10 (O, IN1, IN2);
  output [24:10] O;
  input [14:0] IN1;
  input IN2;
  UB1BPPG_0_10 U0 (O[10], IN1[0], IN2);
  UB1BPPG_1_10 U1 (O[11], IN1[1], IN2);
  UB1BPPG_2_10 U2 (O[12], IN1[2], IN2);
  UB1BPPG_3_10 U3 (O[13], IN1[3], IN2);
  UB1BPPG_4_10 U4 (O[14], IN1[4], IN2);
  UB1BPPG_5_10 U5 (O[15], IN1[5], IN2);
  UB1BPPG_6_10 U6 (O[16], IN1[6], IN2);
  UB1BPPG_7_10 U7 (O[17], IN1[7], IN2);
  UB1BPPG_8_10 U8 (O[18], IN1[8], IN2);
  UB1BPPG_9_10 U9 (O[19], IN1[9], IN2);
  UB1BPPG_10_10 U10 (O[20], IN1[10], IN2);
  UB1BPPG_11_10 U11 (O[21], IN1[11], IN2);
  UB1BPPG_12_10 U12 (O[22], IN1[12], IN2);
  UB1BPPG_13_10 U13 (O[23], IN1[13], IN2);
  UB1BPPG_14_10 U14 (O[24], IN1[14], IN2);
endmodule

module UBVPPG_14_0_12 (O, IN1, IN2);
  output [26:12] O;
  input [14:0] IN1;
  input IN2;
  UB1BPPG_0_12 U0 (O[12], IN1[0], IN2);
  UB1BPPG_1_12 U1 (O[13], IN1[1], IN2);
  UB1BPPG_2_12 U2 (O[14], IN1[2], IN2);
  UB1BPPG_3_12 U3 (O[15], IN1[3], IN2);
  UB1BPPG_4_12 U4 (O[16], IN1[4], IN2);
  UB1BPPG_5_12 U5 (O[17], IN1[5], IN2);
  UB1BPPG_6_12 U6 (O[18], IN1[6], IN2);
  UB1BPPG_7_12 U7 (O[19], IN1[7], IN2);
  UB1BPPG_8_12 U8 (O[20], IN1[8], IN2);
  UB1BPPG_9_12 U9 (O[21], IN1[9], IN2);
  UB1BPPG_10_12 U10 (O[22], IN1[10], IN2);
  UB1BPPG_11_12 U11 (O[23], IN1[11], IN2);
  UB1BPPG_12_12 U12 (O[24], IN1[12], IN2);
  UB1BPPG_13_12 U13 (O[25], IN1[13], IN2);
  UB1BPPG_14_12 U14 (O[26], IN1[14], IN2);
endmodule

module UBVPPG_14_0_14 (O, IN1, IN2);
  output [28:14] O;
  input [14:0] IN1;
  input IN2;
  UB1BPPG_0_14 U0 (O[14], IN1[0], IN2);
  UB1BPPG_1_14 U1 (O[15], IN1[1], IN2);
  UB1BPPG_2_14 U2 (O[16], IN1[2], IN2);
  UB1BPPG_3_14 U3 (O[17], IN1[3], IN2);
  UB1BPPG_4_14 U4 (O[18], IN1[4], IN2);
  UB1BPPG_5_14 U5 (O[19], IN1[5], IN2);
  UB1BPPG_6_14 U6 (O[20], IN1[6], IN2);
  UB1BPPG_7_14 U7 (O[21], IN1[7], IN2);
  UB1BPPG_8_14 U8 (O[22], IN1[8], IN2);
  UB1BPPG_9_14 U9 (O[23], IN1[9], IN2);
  UB1BPPG_10_14 U10 (O[24], IN1[10], IN2);
  UB1BPPG_11_14 U11 (O[25], IN1[11], IN2);
  UB1BPPG_12_14 U12 (O[26], IN1[12], IN2);
  UB1BPPG_13_14 U13 (O[27], IN1[13], IN2);
  UB1BPPG_14_14 U14 (O[28], IN1[14], IN2);
endmodule

module UBVPPG_14_0_2 (O, IN1, IN2);
  output [16:2] O;
  input [14:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
  UB1BPPG_6_2 U6 (O[8], IN1[6], IN2);
  UB1BPPG_7_2 U7 (O[9], IN1[7], IN2);
  UB1BPPG_8_2 U8 (O[10], IN1[8], IN2);
  UB1BPPG_9_2 U9 (O[11], IN1[9], IN2);
  UB1BPPG_10_2 U10 (O[12], IN1[10], IN2);
  UB1BPPG_11_2 U11 (O[13], IN1[11], IN2);
  UB1BPPG_12_2 U12 (O[14], IN1[12], IN2);
  UB1BPPG_13_2 U13 (O[15], IN1[13], IN2);
  UB1BPPG_14_2 U14 (O[16], IN1[14], IN2);
endmodule

module UBVPPG_14_0_4 (O, IN1, IN2);
  output [18:4] O;
  input [14:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
  UB1BPPG_6_4 U6 (O[10], IN1[6], IN2);
  UB1BPPG_7_4 U7 (O[11], IN1[7], IN2);
  UB1BPPG_8_4 U8 (O[12], IN1[8], IN2);
  UB1BPPG_9_4 U9 (O[13], IN1[9], IN2);
  UB1BPPG_10_4 U10 (O[14], IN1[10], IN2);
  UB1BPPG_11_4 U11 (O[15], IN1[11], IN2);
  UB1BPPG_12_4 U12 (O[16], IN1[12], IN2);
  UB1BPPG_13_4 U13 (O[17], IN1[13], IN2);
  UB1BPPG_14_4 U14 (O[18], IN1[14], IN2);
endmodule

module UBVPPG_14_0_6 (O, IN1, IN2);
  output [20:6] O;
  input [14:0] IN1;
  input IN2;
  UB1BPPG_0_6 U0 (O[6], IN1[0], IN2);
  UB1BPPG_1_6 U1 (O[7], IN1[1], IN2);
  UB1BPPG_2_6 U2 (O[8], IN1[2], IN2);
  UB1BPPG_3_6 U3 (O[9], IN1[3], IN2);
  UB1BPPG_4_6 U4 (O[10], IN1[4], IN2);
  UB1BPPG_5_6 U5 (O[11], IN1[5], IN2);
  UB1BPPG_6_6 U6 (O[12], IN1[6], IN2);
  UB1BPPG_7_6 U7 (O[13], IN1[7], IN2);
  UB1BPPG_8_6 U8 (O[14], IN1[8], IN2);
  UB1BPPG_9_6 U9 (O[15], IN1[9], IN2);
  UB1BPPG_10_6 U10 (O[16], IN1[10], IN2);
  UB1BPPG_11_6 U11 (O[17], IN1[11], IN2);
  UB1BPPG_12_6 U12 (O[18], IN1[12], IN2);
  UB1BPPG_13_6 U13 (O[19], IN1[13], IN2);
  UB1BPPG_14_6 U14 (O[20], IN1[14], IN2);
endmodule

module UBVPPG_14_0_8 (O, IN1, IN2);
  output [22:8] O;
  input [14:0] IN1;
  input IN2;
  UB1BPPG_0_8 U0 (O[8], IN1[0], IN2);
  UB1BPPG_1_8 U1 (O[9], IN1[1], IN2);
  UB1BPPG_2_8 U2 (O[10], IN1[2], IN2);
  UB1BPPG_3_8 U3 (O[11], IN1[3], IN2);
  UB1BPPG_4_8 U4 (O[12], IN1[4], IN2);
  UB1BPPG_5_8 U5 (O[13], IN1[5], IN2);
  UB1BPPG_6_8 U6 (O[14], IN1[6], IN2);
  UB1BPPG_7_8 U7 (O[15], IN1[7], IN2);
  UB1BPPG_8_8 U8 (O[16], IN1[8], IN2);
  UB1BPPG_9_8 U9 (O[17], IN1[9], IN2);
  UB1BPPG_10_8 U10 (O[18], IN1[10], IN2);
  UB1BPPG_11_8 U11 (O[19], IN1[11], IN2);
  UB1BPPG_12_8 U12 (O[20], IN1[12], IN2);
  UB1BPPG_13_8 U13 (O[21], IN1[13], IN2);
  UB1BPPG_14_8 U14 (O[22], IN1[14], IN2);
endmodule

