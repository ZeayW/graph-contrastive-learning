/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: Multiplier_5_0_5_000

  Number system: Unsigned binary
  Multiplicand length: 6
  Multiplier length: 6
  Partial product generation: Simple PPG
  Partial product accumulation: Wallace tree
  Final stage addition: Carry-skip adder (variable-block-size)
----------------------------------------------------------------------------*/

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_1(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_2(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_6(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_9(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_10(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBZero_11_11(O);
  output [11:11] O;
  assign O[11] = 0;
endmodule

module UBHA_5(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_5(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_5 U0 (C_0, S_0, X, Y);
  UBHA_5 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_6(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_6 U0 (C_0, S_0, X, Y);
  UBHA_6 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_6_5(Co, S, X, Y, Ci);
  output Co;
  output [6:5] S;
  input Ci;
  input [6:5] X;
  input [6:5] Y;
  wire C6;
  wire C7;
  wire P5;
  wire P6;
  wire Sk;
  assign Sk = ( P5 & P6 ) & Ci;
  assign Co = C7 | Sk;
  UBPFA_5 U0 (C6, S[5], P5, X[5], Y[5], Ci);
  UBPFA_6 U1 (C7, S[6], P6, X[6], Y[6], C6);
endmodule

module UBHA_7(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_7(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_7 U0 (C_0, S_0, X, Y);
  UBHA_7 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_8(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_8(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_8 U0 (C_0, S_0, X, Y);
  UBHA_8 U1 (C_1, S, S_0, Ci);
endmodule

module UBPFA_9(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_9 U0 (C_0, S_0, X, Y);
  UBHA_9 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_9_7(Co, S, X, Y, Ci);
  output Co;
  output [9:7] S;
  input Ci;
  input [9:7] X;
  input [9:7] Y;
  wire C10;
  wire C8;
  wire C9;
  wire P7;
  wire P8;
  wire P9;
  wire Sk;
  assign Sk = ( P7 & P8 & P9 ) & Ci;
  assign Co = C10 | Sk;
  UBPFA_7 U0 (C8, S[7], P7, X[7], Y[7], Ci);
  UBPFA_8 U1 (C9, S[8], P8, X[8], Y[8], C8);
  UBPFA_9 U2 (C10, S[9], P9, X[9], Y[9], C9);
endmodule

module UBPFA_10(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_10 U0 (C_0, S_0, X, Y);
  UBHA_10 U1 (C_1, S, S_0, Ci);
endmodule

module UBHA_11(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBPFA_11(Co, S, P, X, Y, Ci);
  output Co;
  output P;
  output S;
  input Ci;
  input X;
  input Y;
  wire C_0;
  wire C_1;
  wire S_0;
  assign Co = C_0 | C_1;
  assign P = S_0;
  UBHA_11 U0 (C_0, S_0, X, Y);
  UBHA_11 U1 (C_1, S, S_0, Ci);
endmodule

module UBCSkB_11_10(Co, S, X, Y, Ci);
  output Co;
  output [11:10] S;
  input Ci;
  input [11:10] X;
  input [11:10] Y;
  wire C11;
  wire C12;
  wire P10;
  wire P11;
  wire Sk;
  assign Sk = ( P10 & P11 ) & Ci;
  assign Co = C12 | Sk;
  UBPFA_10 U0 (C11, S[10], P10, X[10], Y[10], Ci);
  UBPFA_11 U1 (C12, S[11], P11, X[11], Y[11], C11);
endmodule

module UBPriVCSkA_11_4(S, X, Y, Cin);
  output [12:4] S;
  input Cin;
  input [11:4] X;
  input [11:4] Y;
  wire C10;
  wire C12;
  wire C5;
  wire C7;
  UBFA_4 U0 (C5, S[4], X[4], Y[4], Cin);
  UBCSkB_6_5 U1 (C7, S[6:5], X[6:5], Y[6:5], C5);
  UBCSkB_9_7 U2 (C10, S[9:7], X[9:7], Y[9:7], C7);
  UBCSkB_11_10 U3 (S[12], S[11:10], X[11:10], Y[11:10], C10);
endmodule

module UBZero_4_4(O);
  output [4:4] O;
  assign O[4] = 0;
endmodule

module Multiplier_5_0_5_000(P, IN1, IN2);
  output [11:0] P;
  input [5:0] IN1;
  input [5:0] IN2;
  wire [12:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  MultUB_STD_WAL_VC000 U0 (W, IN1, IN2);
endmodule

module CSA_10_0_8_3_10_5 (C, S, X, Y, Z);
  output [11:4] C;
  output [10:0] S;
  input [10:0] X;
  input [8:3] Y;
  input [10:5] Z;
  UBCON_2_0 U0 (S[2:0], X[2:0]);
  PureCSHA_4_3 U1 (C[5:4], S[4:3], Y[4:3], X[4:3]);
  PureCSA_8_5 U2 (C[9:6], S[8:5], Z[8:5], Y[8:5], X[8:5]);
  PureCSHA_10_9 U3 (C[11:10], S[10:9], Z[10:9], X[10:9]);
endmodule

module CSA_5_0_6_1_7_2 (C, S, X, Y, Z);
  output [7:2] C;
  output [7:0] S;
  input [5:0] X;
  input [6:1] Y;
  input [7:2] Z;
  UB1DCON_0 U0 (S[0], X[0]);
  UBHA_1 U1 (C[2], S[1], Y[1], X[1]);
  PureCSA_5_2 U2 (C[6:3], S[5:2], Z[5:2], Y[5:2], X[5:2]);
  UBHA_6 U3 (C[7], S[6], Z[6], Y[6]);
  UB1DCON_7 U4 (S[7], Z[7]);
endmodule

module CSA_7_0_7_2_10_3 (C, S, X, Y, Z);
  output [8:3] C;
  output [10:0] S;
  input [7:0] X;
  input [7:2] Y;
  input [10:3] Z;
  UBCON_1_0 U0 (S[1:0], X[1:0]);
  UBHA_2 U1 (C[3], S[2], Y[2], X[2]);
  PureCSA_7_3 U2 (C[8:4], S[7:3], Z[7:3], Y[7:3], X[7:3]);
  UBCON_10_8 U3 (S[10:8], Z[10:8]);
endmodule

module CSA_8_3_9_4_10_5 (C, S, X, Y, Z);
  output [10:5] C;
  output [10:3] S;
  input [8:3] X;
  input [9:4] Y;
  input [10:5] Z;
  UB1DCON_3 U0 (S[3], X[3]);
  UBHA_4 U1 (C[5], S[4], Y[4], X[4]);
  PureCSA_8_5 U2 (C[9:6], S[8:5], Z[8:5], Y[8:5], X[8:5]);
  UBHA_9 U3 (C[10], S[9], Z[9], Y[9]);
  UB1DCON_10 U4 (S[10], Z[10]);
endmodule

module MultUB_STD_WAL_VC000 (P, IN1, IN2);
  output [12:0] P;
  input [5:0] IN1;
  input [5:0] IN2;
  wire [5:0] PP0;
  wire [6:1] PP1;
  wire [7:2] PP2;
  wire [8:3] PP3;
  wire [9:4] PP4;
  wire [10:5] PP5;
  wire [11:4] S1;
  wire [10:0] S2;
  UBPPG_5_0_5_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, IN1, IN2);
  WLCTR_5_0_6_1_7_2000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5);
  UBVCSkA_11_4_10_0 U2 (P, S1, S2);
endmodule

module PureCSA_5_2 (C, S, X, Y, Z);
  output [6:3] C;
  output [5:2] S;
  input [5:2] X;
  input [5:2] Y;
  input [5:2] Z;
  UBFA_2 U0 (C[3], S[2], X[2], Y[2], Z[2]);
  UBFA_3 U1 (C[4], S[3], X[3], Y[3], Z[3]);
  UBFA_4 U2 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U3 (C[6], S[5], X[5], Y[5], Z[5]);
endmodule

module PureCSA_7_3 (C, S, X, Y, Z);
  output [8:4] C;
  output [7:3] S;
  input [7:3] X;
  input [7:3] Y;
  input [7:3] Z;
  UBFA_3 U0 (C[4], S[3], X[3], Y[3], Z[3]);
  UBFA_4 U1 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U2 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U3 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U4 (C[8], S[7], X[7], Y[7], Z[7]);
endmodule

module PureCSA_8_5 (C, S, X, Y, Z);
  output [9:6] C;
  output [8:5] S;
  input [8:5] X;
  input [8:5] Y;
  input [8:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U3 (C[9], S[8], X[8], Y[8], Z[8]);
endmodule

module PureCSHA_10_9 (C, S, X, Y);
  output [11:10] C;
  output [10:9] S;
  input [10:9] X;
  input [10:9] Y;
  UBHA_9 U0 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U1 (C[11], S[10], X[10], Y[10]);
endmodule

module PureCSHA_4_3 (C, S, X, Y);
  output [5:4] C;
  output [4:3] S;
  input [4:3] X;
  input [4:3] Y;
  UBHA_3 U0 (C[4], S[3], X[3], Y[3]);
  UBHA_4 U1 (C[5], S[4], X[4], Y[4]);
endmodule

module UBCON_10_4 (O, I);
  output [10:4] O;
  input [10:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
endmodule

module UBCON_10_8 (O, I);
  output [10:8] O;
  input [10:8] I;
  UB1DCON_8 U0 (O[8], I[8]);
  UB1DCON_9 U1 (O[9], I[9]);
  UB1DCON_10 U2 (O[10], I[10]);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBCON_3_0 (O, I);
  output [3:0] O;
  input [3:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
endmodule

module UBExtender_10_4_1000 (O, I);
  output [11:4] O;
  input [10:4] I;
  UBCON_10_4 U0 (O[10:4], I[10:4]);
  UBZero_11_11 U1 (O[11]);
endmodule

module UBPPG_5_0_5_0 (PP0, PP1, PP2, PP3, PP4, PP5, IN1, IN2);
  output [5:0] PP0;
  output [6:1] PP1;
  output [7:2] PP2;
  output [8:3] PP3;
  output [9:4] PP4;
  output [10:5] PP5;
  input [5:0] IN1;
  input [5:0] IN2;
  UBVPPG_5_0_0 U0 (PP0, IN1, IN2[0]);
  UBVPPG_5_0_1 U1 (PP1, IN1, IN2[1]);
  UBVPPG_5_0_2 U2 (PP2, IN1, IN2[2]);
  UBVPPG_5_0_3 U3 (PP3, IN1, IN2[3]);
  UBVPPG_5_0_4 U4 (PP4, IN1, IN2[4]);
  UBVPPG_5_0_5 U5 (PP5, IN1, IN2[5]);
endmodule

module UBPureVCSkA_11_4 (S, X, Y);
  output [12:4] S;
  input [11:4] X;
  input [11:4] Y;
  wire C;
  UBPriVCSkA_11_4 U0 (S, X, Y, C);
  UBZero_4_4 U1 (C);
endmodule

module UBVCSkA_11_4_10_0 (S, X, Y);
  output [12:0] S;
  input [11:4] X;
  input [10:0] Y;
  wire [11:4] Z;
  UBExtender_10_4_1000 U0 (Z[11:4], Y[10:4]);
  UBPureVCSkA_11_4 U1 (S[12:4], X[11:4], Z[11:4]);
  UBCON_3_0 U2 (S[3:0], Y[3:0]);
endmodule

module UBVPPG_5_0_0 (O, IN1, IN2);
  output [5:0] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
endmodule

module UBVPPG_5_0_1 (O, IN1, IN2);
  output [6:1] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_1 U0 (O[1], IN1[0], IN2);
  UB1BPPG_1_1 U1 (O[2], IN1[1], IN2);
  UB1BPPG_2_1 U2 (O[3], IN1[2], IN2);
  UB1BPPG_3_1 U3 (O[4], IN1[3], IN2);
  UB1BPPG_4_1 U4 (O[5], IN1[4], IN2);
  UB1BPPG_5_1 U5 (O[6], IN1[5], IN2);
endmodule

module UBVPPG_5_0_2 (O, IN1, IN2);
  output [7:2] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
endmodule

module UBVPPG_5_0_3 (O, IN1, IN2);
  output [8:3] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_3 U0 (O[3], IN1[0], IN2);
  UB1BPPG_1_3 U1 (O[4], IN1[1], IN2);
  UB1BPPG_2_3 U2 (O[5], IN1[2], IN2);
  UB1BPPG_3_3 U3 (O[6], IN1[3], IN2);
  UB1BPPG_4_3 U4 (O[7], IN1[4], IN2);
  UB1BPPG_5_3 U5 (O[8], IN1[5], IN2);
endmodule

module UBVPPG_5_0_4 (O, IN1, IN2);
  output [9:4] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
endmodule

module UBVPPG_5_0_5 (O, IN1, IN2);
  output [10:5] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_5 U0 (O[5], IN1[0], IN2);
  UB1BPPG_1_5 U1 (O[6], IN1[1], IN2);
  UB1BPPG_2_5 U2 (O[7], IN1[2], IN2);
  UB1BPPG_3_5 U3 (O[8], IN1[3], IN2);
  UB1BPPG_4_5 U4 (O[9], IN1[4], IN2);
  UB1BPPG_5_5 U5 (O[10], IN1[5], IN2);
endmodule

module WLCTR_5_0_6_1_7_2000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5);
  output [11:4] S1;
  output [10:0] S2;
  input [5:0] PP0;
  input [6:1] PP1;
  input [7:2] PP2;
  input [8:3] PP3;
  input [9:4] PP4;
  input [10:5] PP5;
  wire [7:2] IC0;
  wire [10:5] IC1;
  wire [8:3] IC2;
  wire [7:0] IS0;
  wire [10:3] IS1;
  wire [10:0] IS2;
  CSA_5_0_6_1_7_2 U0 (IC0, IS0, PP0, PP1, PP2);
  CSA_8_3_9_4_10_5 U1 (IC1, IS1, PP3, PP4, PP5);
  CSA_7_0_7_2_10_3 U2 (IC2, IS2, IS0, IC0, IS1);
  CSA_10_0_8_3_10_5 U3 (S1, S2, IS2, IC2, IC1);
endmodule

