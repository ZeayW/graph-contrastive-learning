/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: Multiplier_5_0_5_000

  Number system: Unsigned binary
  Multiplicand length: 6
  Multiplier length: 6
  Partial product generation: Simple PPG
  Partial product accumulation: Balanced delay tree
  Final stage addition: Ripple carry adder
----------------------------------------------------------------------------*/

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_1(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_2(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_6(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_9(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_8(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_10(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBZero_3_3(O);
  output [3:3] O;
  assign O[3] = 0;
endmodule

module Multiplier_5_0_5_000(P, IN1, IN2);
  output [11:0] P;
  input [5:0] IN1;
  input [5:0] IN2;
  wire [12:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  MultUB_STD_BLD_RC000 U0 (W, IN1, IN2);
endmodule

module BLDCON_7_2_7_0_10000 (S1, S2, IN0, IN1, IN2, IN3);
  output [11:3] S1;
  output [11:0] S2;
  input [7:2] IN0;
  input [7:0] IN1;
  input [10:5] IN2;
  input [10:3] IN3;
  wire [11:4] W1;
  wire [10:0] W2;
  CSA_7_0_10_5_10_3 U0 (W1, W2, IN1, IN2, IN3);
  CSA_11_4_10_0_7_2 U1 (S1, S2, W1, W2, IN0);
endmodule

module BLDTR_5_0_6_1_7_2000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5);
  output [11:3] S1;
  output [11:0] S2;
  input [5:0] PP0;
  input [6:1] PP1;
  input [7:2] PP2;
  input [8:3] PP3;
  input [9:4] PP4;
  input [10:5] PP5;
  wire [7:2] W0;
  wire [7:0] W1;
  wire [10:5] W2;
  wire [10:3] W3;
  UBARYACC_5_0_6_1_000 U0 (W0, W1, PP0, PP1, PP2);
  UBARYACC_8_3_9_4_000 U1 (W2, W3, PP3, PP4, PP5);
  BLDCON_7_2_7_0_10000 U2 (S1, S2, W0, W1, W2, W3);
endmodule

module CSA_11_4_10_0_7_2 (C, S, X, Y, Z);
  output [11:3] C;
  output [11:0] S;
  input [11:4] X;
  input [10:0] Y;
  input [7:2] Z;
  UBCON_1_0 U0 (S[1:0], Y[1:0]);
  PureCSHA_3_2 U1 (C[4:3], S[3:2], Z[3:2], Y[3:2]);
  PureCSA_7_4 U2 (C[8:5], S[7:4], X[7:4], Z[7:4], Y[7:4]);
  PureCSHA_10_8 U3 (C[11:9], S[10:8], X[10:8], Y[10:8]);
  UB1DCON_11 U4 (S[11], X[11]);
endmodule

module CSA_5_0_6_1_7_2 (C, S, X, Y, Z);
  output [7:2] C;
  output [7:0] S;
  input [5:0] X;
  input [6:1] Y;
  input [7:2] Z;
  UB1DCON_0 U0 (S[0], X[0]);
  UBHA_1 U1 (C[2], S[1], Y[1], X[1]);
  PureCSA_5_2 U2 (C[6:3], S[5:2], Z[5:2], Y[5:2], X[5:2]);
  UBHA_6 U3 (C[7], S[6], Z[6], Y[6]);
  UB1DCON_7 U4 (S[7], Z[7]);
endmodule

module CSA_7_0_10_5_10_3 (C, S, X, Y, Z);
  output [11:4] C;
  output [10:0] S;
  input [7:0] X;
  input [10:5] Y;
  input [10:3] Z;
  UBCON_2_0 U0 (S[2:0], X[2:0]);
  PureCSHA_4_3 U1 (C[5:4], S[4:3], Z[4:3], X[4:3]);
  PureCSA_7_5 U2 (C[8:6], S[7:5], Y[7:5], Z[7:5], X[7:5]);
  PureCSHA_10_8 U3 (C[11:9], S[10:8], Z[10:8], Y[10:8]);
endmodule

module CSA_8_3_9_4_10_5 (C, S, X, Y, Z);
  output [10:5] C;
  output [10:3] S;
  input [8:3] X;
  input [9:4] Y;
  input [10:5] Z;
  UB1DCON_3 U0 (S[3], X[3]);
  UBHA_4 U1 (C[5], S[4], Y[4], X[4]);
  PureCSA_8_5 U2 (C[9:6], S[8:5], Z[8:5], Y[8:5], X[8:5]);
  UBHA_9 U3 (C[10], S[9], Z[9], Y[9]);
  UB1DCON_10 U4 (S[10], Z[10]);
endmodule

module MultUB_STD_BLD_RC000 (P, IN1, IN2);
  output [12:0] P;
  input [5:0] IN1;
  input [5:0] IN2;
  wire [5:0] PP0;
  wire [6:1] PP1;
  wire [7:2] PP2;
  wire [8:3] PP3;
  wire [9:4] PP4;
  wire [10:5] PP5;
  wire [11:3] S1;
  wire [11:0] S2;
  UBPPG_5_0_5_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, IN1, IN2);
  BLDTR_5_0_6_1_7_2000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5);
  UBRCA_11_3_11_0 U2 (P, S1, S2);
endmodule

module PureCSA_5_2 (C, S, X, Y, Z);
  output [6:3] C;
  output [5:2] S;
  input [5:2] X;
  input [5:2] Y;
  input [5:2] Z;
  UBFA_2 U0 (C[3], S[2], X[2], Y[2], Z[2]);
  UBFA_3 U1 (C[4], S[3], X[3], Y[3], Z[3]);
  UBFA_4 U2 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U3 (C[6], S[5], X[5], Y[5], Z[5]);
endmodule

module PureCSA_7_4 (C, S, X, Y, Z);
  output [8:5] C;
  output [7:4] S;
  input [7:4] X;
  input [7:4] Y;
  input [7:4] Z;
  UBFA_4 U0 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U1 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U2 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U3 (C[8], S[7], X[7], Y[7], Z[7]);
endmodule

module PureCSA_7_5 (C, S, X, Y, Z);
  output [8:6] C;
  output [7:5] S;
  input [7:5] X;
  input [7:5] Y;
  input [7:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
endmodule

module PureCSA_8_5 (C, S, X, Y, Z);
  output [9:6] C;
  output [8:5] S;
  input [8:5] X;
  input [8:5] Y;
  input [8:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U3 (C[9], S[8], X[8], Y[8], Z[8]);
endmodule

module PureCSHA_10_8 (C, S, X, Y);
  output [11:9] C;
  output [10:8] S;
  input [10:8] X;
  input [10:8] Y;
  UBHA_8 U0 (C[9], S[8], X[8], Y[8]);
  UBHA_9 U1 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U2 (C[11], S[10], X[10], Y[10]);
endmodule

module PureCSHA_3_2 (C, S, X, Y);
  output [4:3] C;
  output [3:2] S;
  input [3:2] X;
  input [3:2] Y;
  UBHA_2 U0 (C[3], S[2], X[2], Y[2]);
  UBHA_3 U1 (C[4], S[3], X[3], Y[3]);
endmodule

module PureCSHA_4_3 (C, S, X, Y);
  output [5:4] C;
  output [4:3] S;
  input [4:3] X;
  input [4:3] Y;
  UBHA_3 U0 (C[4], S[3], X[3], Y[3]);
  UBHA_4 U1 (C[5], S[4], X[4], Y[4]);
endmodule

module UBARYACC_5_0_6_1_000 (S1, S2, PP0, PP1, PP2);
  output [7:2] S1;
  output [7:0] S2;
  input [5:0] PP0;
  input [6:1] PP1;
  input [7:2] PP2;
  CSA_5_0_6_1_7_2 U0 (S1, S2, PP0, PP1, PP2);
endmodule

module UBARYACC_8_3_9_4_000 (S1, S2, PP0, PP1, PP2);
  output [10:5] S1;
  output [10:3] S2;
  input [8:3] PP0;
  input [9:4] PP1;
  input [10:5] PP2;
  CSA_8_3_9_4_10_5 U0 (S1, S2, PP0, PP1, PP2);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBPPG_5_0_5_0 (PP0, PP1, PP2, PP3, PP4, PP5, IN1, IN2);
  output [5:0] PP0;
  output [6:1] PP1;
  output [7:2] PP2;
  output [8:3] PP3;
  output [9:4] PP4;
  output [10:5] PP5;
  input [5:0] IN1;
  input [5:0] IN2;
  UBVPPG_5_0_0 U0 (PP0, IN1, IN2[0]);
  UBVPPG_5_0_1 U1 (PP1, IN1, IN2[1]);
  UBVPPG_5_0_2 U2 (PP2, IN1, IN2[2]);
  UBVPPG_5_0_3 U3 (PP3, IN1, IN2[3]);
  UBVPPG_5_0_4 U4 (PP4, IN1, IN2[4]);
  UBVPPG_5_0_5 U5 (PP5, IN1, IN2[5]);
endmodule

module UBPriRCA_11_3 (S, X, Y, Cin);
  output [12:3] S;
  input Cin;
  input [11:3] X;
  input [11:3] Y;
  wire C10;
  wire C11;
  wire C4;
  wire C5;
  wire C6;
  wire C7;
  wire C8;
  wire C9;
  UBFA_3 U0 (C4, S[3], X[3], Y[3], Cin);
  UBFA_4 U1 (C5, S[4], X[4], Y[4], C4);
  UBFA_5 U2 (C6, S[5], X[5], Y[5], C5);
  UBFA_6 U3 (C7, S[6], X[6], Y[6], C6);
  UBFA_7 U4 (C8, S[7], X[7], Y[7], C7);
  UBFA_8 U5 (C9, S[8], X[8], Y[8], C8);
  UBFA_9 U6 (C10, S[9], X[9], Y[9], C9);
  UBFA_10 U7 (C11, S[10], X[10], Y[10], C10);
  UBFA_11 U8 (S[12], S[11], X[11], Y[11], C11);
endmodule

module UBPureRCA_11_3 (S, X, Y);
  output [12:3] S;
  input [11:3] X;
  input [11:3] Y;
  wire C;
  UBPriRCA_11_3 U0 (S, X, Y, C);
  UBZero_3_3 U1 (C);
endmodule

module UBRCA_11_3_11_0 (S, X, Y);
  output [12:0] S;
  input [11:3] X;
  input [11:0] Y;
  UBPureRCA_11_3 U0 (S[12:3], X[11:3], Y[11:3]);
  UBCON_2_0 U1 (S[2:0], Y[2:0]);
endmodule

module UBVPPG_5_0_0 (O, IN1, IN2);
  output [5:0] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
endmodule

module UBVPPG_5_0_1 (O, IN1, IN2);
  output [6:1] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_1 U0 (O[1], IN1[0], IN2);
  UB1BPPG_1_1 U1 (O[2], IN1[1], IN2);
  UB1BPPG_2_1 U2 (O[3], IN1[2], IN2);
  UB1BPPG_3_1 U3 (O[4], IN1[3], IN2);
  UB1BPPG_4_1 U4 (O[5], IN1[4], IN2);
  UB1BPPG_5_1 U5 (O[6], IN1[5], IN2);
endmodule

module UBVPPG_5_0_2 (O, IN1, IN2);
  output [7:2] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
endmodule

module UBVPPG_5_0_3 (O, IN1, IN2);
  output [8:3] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_3 U0 (O[3], IN1[0], IN2);
  UB1BPPG_1_3 U1 (O[4], IN1[1], IN2);
  UB1BPPG_2_3 U2 (O[5], IN1[2], IN2);
  UB1BPPG_3_3 U3 (O[6], IN1[3], IN2);
  UB1BPPG_4_3 U4 (O[7], IN1[4], IN2);
  UB1BPPG_5_3 U5 (O[8], IN1[5], IN2);
endmodule

module UBVPPG_5_0_4 (O, IN1, IN2);
  output [9:4] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
endmodule

module UBVPPG_5_0_5 (O, IN1, IN2);
  output [10:5] O;
  input [5:0] IN1;
  input IN2;
  UB1BPPG_0_5 U0 (O[5], IN1[0], IN2);
  UB1BPPG_1_5 U1 (O[6], IN1[1], IN2);
  UB1BPPG_2_5 U2 (O[7], IN1[2], IN2);
  UB1BPPG_3_5 U3 (O[8], IN1[3], IN2);
  UB1BPPG_4_5 U4 (O[9], IN1[4], IN2);
  UB1BPPG_5_5 U5 (O[10], IN1[5], IN2);
endmodule

