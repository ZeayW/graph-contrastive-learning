library IEEE;
use IEEE.std_logic_1164.all;
entity CSA_10_0_10_3_11_000 is
  port(
      C : out std_logic_vector(11 downto 4);
      S : out std_logic_vector(11 downto 0);
      X : in std_logic_vector(10 downto 0);
      Y : in std_logic_vector(10 downto 3);
      Z : in std_logic_vector(11 downto 4));
end CSA_10_0_10_3_11_000;

architecture CSA_10_0_10_3_11_000 of CSA_10_0_10_3_11_000 is
  component UBCON_2_0 
    port(
      O : out std_logic_vector(2 downto 0);
      I : in std_logic_vector(2 downto 0));
  end component;
  component UBHA_3 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic);
  end component;
  component PureCSA_10_4 
    port(
      C : out std_logic_vector(11 downto 5);
      S : out std_logic_vector(10 downto 4);
      X : in std_logic_vector(10 downto 4);
      Y : in std_logic_vector(10 downto 4);
      Z : in std_logic_vector(10 downto 4));
  end component;
  component UB1DCON_11 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
begin
  U0: UBCON_2_0 port map (S(2 downto 0), X(2 downto 0));
  U1: UBHA_3 port map (C(4), S(3), Y(3), X(3));
  U2: PureCSA_10_4 port map (C(11 downto 5), S(10 downto 4), Z(10 downto 4), Y(10 downto 4), X(10 downto 4));
  U3: UB1DCON_11 port map (S(11), Z(11));
end CSA_10_0_10_3_11_000;

library IEEE;
use IEEE.std_logic_1164.all;
entity CSA_11_0_11_4_12_000 is
  port(
      C : out std_logic_vector(12 downto 5);
      S : out std_logic_vector(12 downto 0);
      X : in std_logic_vector(11 downto 0);
      Y : in std_logic_vector(11 downto 4);
      Z : in std_logic_vector(12 downto 5));
end CSA_11_0_11_4_12_000;

architecture CSA_11_0_11_4_12_000 of CSA_11_0_11_4_12_000 is
  component UBCON_3_0 
    port(
      O : out std_logic_vector(3 downto 0);
      I : in std_logic_vector(3 downto 0));
  end component;
  component UBHA_4 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic);
  end component;
  component PureCSA_11_5 
    port(
      C : out std_logic_vector(12 downto 6);
      S : out std_logic_vector(11 downto 5);
      X : in std_logic_vector(11 downto 5);
      Y : in std_logic_vector(11 downto 5);
      Z : in std_logic_vector(11 downto 5));
  end component;
  component UB1DCON_12 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
begin
  U0: UBCON_3_0 port map (S(3 downto 0), X(3 downto 0));
  U1: UBHA_4 port map (C(5), S(4), Y(4), X(4));
  U2: PureCSA_11_5 port map (C(12 downto 6), S(11 downto 5), Z(11 downto 5), Y(11 downto 5), X(11 downto 5));
  U3: UB1DCON_12 port map (S(12), Z(12));
end CSA_11_0_11_4_12_000;

library IEEE;
use IEEE.std_logic_1164.all;
entity CSA_12_0_12_5_13_000 is
  port(
      C : out std_logic_vector(13 downto 6);
      S : out std_logic_vector(13 downto 0);
      X : in std_logic_vector(12 downto 0);
      Y : in std_logic_vector(12 downto 5);
      Z : in std_logic_vector(13 downto 6));
end CSA_12_0_12_5_13_000;

architecture CSA_12_0_12_5_13_000 of CSA_12_0_12_5_13_000 is
  component UBCON_4_0 
    port(
      O : out std_logic_vector(4 downto 0);
      I : in std_logic_vector(4 downto 0));
  end component;
  component UBHA_5 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic);
  end component;
  component PureCSA_12_6 
    port(
      C : out std_logic_vector(13 downto 7);
      S : out std_logic_vector(12 downto 6);
      X : in std_logic_vector(12 downto 6);
      Y : in std_logic_vector(12 downto 6);
      Z : in std_logic_vector(12 downto 6));
  end component;
  component UB1DCON_13 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
begin
  U0: UBCON_4_0 port map (S(4 downto 0), X(4 downto 0));
  U1: UBHA_5 port map (C(6), S(5), Y(5), X(5));
  U2: PureCSA_12_6 port map (C(13 downto 7), S(12 downto 6), Z(12 downto 6), Y(12 downto 6), X(12 downto 6));
  U3: UB1DCON_13 port map (S(13), Z(13));
end CSA_12_0_12_5_13_000;

library IEEE;
use IEEE.std_logic_1164.all;
entity CSA_13_0_13_6_14_000 is
  port(
      C : out std_logic_vector(14 downto 7);
      S : out std_logic_vector(14 downto 0);
      X : in std_logic_vector(13 downto 0);
      Y : in std_logic_vector(13 downto 6);
      Z : in std_logic_vector(14 downto 7));
end CSA_13_0_13_6_14_000;

architecture CSA_13_0_13_6_14_000 of CSA_13_0_13_6_14_000 is
  component UBCON_5_0 
    port(
      O : out std_logic_vector(5 downto 0);
      I : in std_logic_vector(5 downto 0));
  end component;
  component UBHA_6 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic);
  end component;
  component PureCSA_13_7 
    port(
      C : out std_logic_vector(14 downto 8);
      S : out std_logic_vector(13 downto 7);
      X : in std_logic_vector(13 downto 7);
      Y : in std_logic_vector(13 downto 7);
      Z : in std_logic_vector(13 downto 7));
  end component;
  component UB1DCON_14 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
begin
  U0: UBCON_5_0 port map (S(5 downto 0), X(5 downto 0));
  U1: UBHA_6 port map (C(7), S(6), Y(6), X(6));
  U2: PureCSA_13_7 port map (C(14 downto 8), S(13 downto 7), Z(13 downto 7), Y(13 downto 7), X(13 downto 7));
  U3: UB1DCON_14 port map (S(14), Z(14));
end CSA_13_0_13_6_14_000;

library IEEE;
use IEEE.std_logic_1164.all;
entity CSA_7_0_8_1_9_2 is
  port(
      C : out std_logic_vector(9 downto 2);
      S : out std_logic_vector(9 downto 0);
      X : in std_logic_vector(7 downto 0);
      Y : in std_logic_vector(8 downto 1);
      Z : in std_logic_vector(9 downto 2));
end CSA_7_0_8_1_9_2;

architecture CSA_7_0_8_1_9_2 of CSA_7_0_8_1_9_2 is
  component UB1DCON_0 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UBHA_1 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic);
  end component;
  component PureCSA_7_2 
    port(
      C : out std_logic_vector(8 downto 3);
      S : out std_logic_vector(7 downto 2);
      X : in std_logic_vector(7 downto 2);
      Y : in std_logic_vector(7 downto 2);
      Z : in std_logic_vector(7 downto 2));
  end component;
  component UBHA_8 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic);
  end component;
  component UB1DCON_9 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
begin
  U0: UB1DCON_0 port map (S(0), X(0));
  U1: UBHA_1 port map (C(2), S(1), Y(1), X(1));
  U2: PureCSA_7_2 port map (C(8 downto 3), S(7 downto 2), Z(7 downto 2), Y(7 downto 2), X(7 downto 2));
  U3: UBHA_8 port map (C(9), S(8), Z(8), Y(8));
  U4: UB1DCON_9 port map (S(9), Z(9));
end CSA_7_0_8_1_9_2;

library IEEE;
use IEEE.std_logic_1164.all;
entity CSA_9_0_9_2_10_3 is
  port(
      C : out std_logic_vector(10 downto 3);
      S : out std_logic_vector(10 downto 0);
      X : in std_logic_vector(9 downto 0);
      Y : in std_logic_vector(9 downto 2);
      Z : in std_logic_vector(10 downto 3));
end CSA_9_0_9_2_10_3;

architecture CSA_9_0_9_2_10_3 of CSA_9_0_9_2_10_3 is
  component UBCON_1_0 
    port(
      O : out std_logic_vector(1 downto 0);
      I : in std_logic_vector(1 downto 0));
  end component;
  component UBHA_2 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic);
  end component;
  component PureCSA_9_3 
    port(
      C : out std_logic_vector(10 downto 4);
      S : out std_logic_vector(9 downto 3);
      X : in std_logic_vector(9 downto 3);
      Y : in std_logic_vector(9 downto 3);
      Z : in std_logic_vector(9 downto 3));
  end component;
  component UB1DCON_10 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
begin
  U0: UBCON_1_0 port map (S(1 downto 0), X(1 downto 0));
  U1: UBHA_2 port map (C(3), S(2), Y(2), X(2));
  U2: PureCSA_9_3 port map (C(10 downto 4), S(9 downto 3), Z(9 downto 3), Y(9 downto 3), X(9 downto 3));
  U3: UB1DCON_10 port map (S(10), Z(10));
end CSA_9_0_9_2_10_3;

library IEEE;
use IEEE.std_logic_1164.all;
entity MultUB_STD_ARY_HC000 is
  port(
      P : out std_logic_vector(15 downto 0);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic_vector(7 downto 0));
end MultUB_STD_ARY_HC000;

architecture MultUB_STD_ARY_HC000 of MultUB_STD_ARY_HC000 is
  component UBPPG_7_0_7_0 
    port(
      PP0 : out std_logic_vector(7 downto 0);
      PP1 : out std_logic_vector(8 downto 1);
      PP2 : out std_logic_vector(9 downto 2);
      PP3 : out std_logic_vector(10 downto 3);
      PP4 : out std_logic_vector(11 downto 4);
      PP5 : out std_logic_vector(12 downto 5);
      PP6 : out std_logic_vector(13 downto 6);
      PP7 : out std_logic_vector(14 downto 7);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic_vector(7 downto 0));
  end component;
  component UBARYACC_7_0_8_1_000 
    port(
      S1 : out std_logic_vector(14 downto 7);
      S2 : out std_logic_vector(14 downto 0);
      PP0 : in std_logic_vector(7 downto 0);
      PP1 : in std_logic_vector(8 downto 1);
      PP2 : in std_logic_vector(9 downto 2);
      PP3 : in std_logic_vector(10 downto 3);
      PP4 : in std_logic_vector(11 downto 4);
      PP5 : in std_logic_vector(12 downto 5);
      PP6 : in std_logic_vector(13 downto 6);
      PP7 : in std_logic_vector(14 downto 7));
  end component;
  component UBHCA_14_7_14_0 
    port(
      S : out std_logic_vector(15 downto 0);
      X : in std_logic_vector(14 downto 7);
      Y : in std_logic_vector(14 downto 0));
  end component;
  signal PP0 : std_logic_vector(7 downto 0);
  signal PP1 : std_logic_vector(8 downto 1);
  signal PP2 : std_logic_vector(9 downto 2);
  signal PP3 : std_logic_vector(10 downto 3);
  signal PP4 : std_logic_vector(11 downto 4);
  signal PP5 : std_logic_vector(12 downto 5);
  signal PP6 : std_logic_vector(13 downto 6);
  signal PP7 : std_logic_vector(14 downto 7);
  signal S1 : std_logic_vector(14 downto 7);
  signal S2 : std_logic_vector(14 downto 0);
begin
  U0: UBPPG_7_0_7_0 port map (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, IN1, IN2);
  U1: UBARYACC_7_0_8_1_000 port map (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7);
  U2: UBHCA_14_7_14_0 port map (P, S1, S2);
end MultUB_STD_ARY_HC000;

library IEEE;
use IEEE.std_logic_1164.all;
entity PureCSA_10_4 is
  port(
      C : out std_logic_vector(11 downto 5);
      S : out std_logic_vector(10 downto 4);
      X : in std_logic_vector(10 downto 4);
      Y : in std_logic_vector(10 downto 4);
      Z : in std_logic_vector(10 downto 4));
end PureCSA_10_4;

architecture PureCSA_10_4 of PureCSA_10_4 is
  component UBFA_4 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_5 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_6 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_7 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_8 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_9 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_10 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
begin
  U0: UBFA_4 port map (C(5), S(4), X(4), Y(4), Z(4));
  U1: UBFA_5 port map (C(6), S(5), X(5), Y(5), Z(5));
  U2: UBFA_6 port map (C(7), S(6), X(6), Y(6), Z(6));
  U3: UBFA_7 port map (C(8), S(7), X(7), Y(7), Z(7));
  U4: UBFA_8 port map (C(9), S(8), X(8), Y(8), Z(8));
  U5: UBFA_9 port map (C(10), S(9), X(9), Y(9), Z(9));
  U6: UBFA_10 port map (C(11), S(10), X(10), Y(10), Z(10));
end PureCSA_10_4;

library IEEE;
use IEEE.std_logic_1164.all;
entity PureCSA_11_5 is
  port(
      C : out std_logic_vector(12 downto 6);
      S : out std_logic_vector(11 downto 5);
      X : in std_logic_vector(11 downto 5);
      Y : in std_logic_vector(11 downto 5);
      Z : in std_logic_vector(11 downto 5));
end PureCSA_11_5;

architecture PureCSA_11_5 of PureCSA_11_5 is
  component UBFA_5 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_6 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_7 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_8 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_9 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_10 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_11 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
begin
  U0: UBFA_5 port map (C(6), S(5), X(5), Y(5), Z(5));
  U1: UBFA_6 port map (C(7), S(6), X(6), Y(6), Z(6));
  U2: UBFA_7 port map (C(8), S(7), X(7), Y(7), Z(7));
  U3: UBFA_8 port map (C(9), S(8), X(8), Y(8), Z(8));
  U4: UBFA_9 port map (C(10), S(9), X(9), Y(9), Z(9));
  U5: UBFA_10 port map (C(11), S(10), X(10), Y(10), Z(10));
  U6: UBFA_11 port map (C(12), S(11), X(11), Y(11), Z(11));
end PureCSA_11_5;

library IEEE;
use IEEE.std_logic_1164.all;
entity PureCSA_12_6 is
  port(
      C : out std_logic_vector(13 downto 7);
      S : out std_logic_vector(12 downto 6);
      X : in std_logic_vector(12 downto 6);
      Y : in std_logic_vector(12 downto 6);
      Z : in std_logic_vector(12 downto 6));
end PureCSA_12_6;

architecture PureCSA_12_6 of PureCSA_12_6 is
  component UBFA_6 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_7 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_8 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_9 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_10 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_11 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_12 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
begin
  U0: UBFA_6 port map (C(7), S(6), X(6), Y(6), Z(6));
  U1: UBFA_7 port map (C(8), S(7), X(7), Y(7), Z(7));
  U2: UBFA_8 port map (C(9), S(8), X(8), Y(8), Z(8));
  U3: UBFA_9 port map (C(10), S(9), X(9), Y(9), Z(9));
  U4: UBFA_10 port map (C(11), S(10), X(10), Y(10), Z(10));
  U5: UBFA_11 port map (C(12), S(11), X(11), Y(11), Z(11));
  U6: UBFA_12 port map (C(13), S(12), X(12), Y(12), Z(12));
end PureCSA_12_6;

library IEEE;
use IEEE.std_logic_1164.all;
entity PureCSA_13_7 is
  port(
      C : out std_logic_vector(14 downto 8);
      S : out std_logic_vector(13 downto 7);
      X : in std_logic_vector(13 downto 7);
      Y : in std_logic_vector(13 downto 7);
      Z : in std_logic_vector(13 downto 7));
end PureCSA_13_7;

architecture PureCSA_13_7 of PureCSA_13_7 is
  component UBFA_7 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_8 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_9 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_10 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_11 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_12 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_13 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
begin
  U0: UBFA_7 port map (C(8), S(7), X(7), Y(7), Z(7));
  U1: UBFA_8 port map (C(9), S(8), X(8), Y(8), Z(8));
  U2: UBFA_9 port map (C(10), S(9), X(9), Y(9), Z(9));
  U3: UBFA_10 port map (C(11), S(10), X(10), Y(10), Z(10));
  U4: UBFA_11 port map (C(12), S(11), X(11), Y(11), Z(11));
  U5: UBFA_12 port map (C(13), S(12), X(12), Y(12), Z(12));
  U6: UBFA_13 port map (C(14), S(13), X(13), Y(13), Z(13));
end PureCSA_13_7;

library IEEE;
use IEEE.std_logic_1164.all;
entity PureCSA_7_2 is
  port(
      C : out std_logic_vector(8 downto 3);
      S : out std_logic_vector(7 downto 2);
      X : in std_logic_vector(7 downto 2);
      Y : in std_logic_vector(7 downto 2);
      Z : in std_logic_vector(7 downto 2));
end PureCSA_7_2;

architecture PureCSA_7_2 of PureCSA_7_2 is
  component UBFA_2 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_3 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_4 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_5 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_6 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_7 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
begin
  U0: UBFA_2 port map (C(3), S(2), X(2), Y(2), Z(2));
  U1: UBFA_3 port map (C(4), S(3), X(3), Y(3), Z(3));
  U2: UBFA_4 port map (C(5), S(4), X(4), Y(4), Z(4));
  U3: UBFA_5 port map (C(6), S(5), X(5), Y(5), Z(5));
  U4: UBFA_6 port map (C(7), S(6), X(6), Y(6), Z(6));
  U5: UBFA_7 port map (C(8), S(7), X(7), Y(7), Z(7));
end PureCSA_7_2;

library IEEE;
use IEEE.std_logic_1164.all;
entity PureCSA_9_3 is
  port(
      C : out std_logic_vector(10 downto 4);
      S : out std_logic_vector(9 downto 3);
      X : in std_logic_vector(9 downto 3);
      Y : in std_logic_vector(9 downto 3);
      Z : in std_logic_vector(9 downto 3));
end PureCSA_9_3;

architecture PureCSA_9_3 of PureCSA_9_3 is
  component UBFA_3 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_4 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_5 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_6 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_7 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_8 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
  component UBFA_9 
    port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
  end component;
begin
  U0: UBFA_3 port map (C(4), S(3), X(3), Y(3), Z(3));
  U1: UBFA_4 port map (C(5), S(4), X(4), Y(4), Z(4));
  U2: UBFA_5 port map (C(6), S(5), X(5), Y(5), Z(5));
  U3: UBFA_6 port map (C(7), S(6), X(6), Y(6), Z(6));
  U4: UBFA_7 port map (C(8), S(7), X(7), Y(7), Z(7));
  U5: UBFA_8 port map (C(9), S(8), X(8), Y(8), Z(8));
  U6: UBFA_9 port map (C(10), S(9), X(9), Y(9), Z(9));
end PureCSA_9_3;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_0_0 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_0_0;

architecture UB1BPPG_0_0 of UB1BPPG_0_0 is
begin
-- TODO
end UB1BPPG_0_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_0_1 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_0_1;

architecture UB1BPPG_0_1 of UB1BPPG_0_1 is
begin
-- TODO
end UB1BPPG_0_1;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_0_2 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_0_2;

architecture UB1BPPG_0_2 of UB1BPPG_0_2 is
begin
-- TODO
end UB1BPPG_0_2;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_0_3 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_0_3;

architecture UB1BPPG_0_3 of UB1BPPG_0_3 is
begin
-- TODO
end UB1BPPG_0_3;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_0_4 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_0_4;

architecture UB1BPPG_0_4 of UB1BPPG_0_4 is
begin
-- TODO
end UB1BPPG_0_4;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_0_5 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_0_5;

architecture UB1BPPG_0_5 of UB1BPPG_0_5 is
begin
-- TODO
end UB1BPPG_0_5;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_0_6 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_0_6;

architecture UB1BPPG_0_6 of UB1BPPG_0_6 is
begin
-- TODO
end UB1BPPG_0_6;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_0_7 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_0_7;

architecture UB1BPPG_0_7 of UB1BPPG_0_7 is
begin
-- TODO
end UB1BPPG_0_7;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_1_0 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_1_0;

architecture UB1BPPG_1_0 of UB1BPPG_1_0 is
begin
-- TODO
end UB1BPPG_1_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_1_1 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_1_1;

architecture UB1BPPG_1_1 of UB1BPPG_1_1 is
begin
-- TODO
end UB1BPPG_1_1;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_1_2 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_1_2;

architecture UB1BPPG_1_2 of UB1BPPG_1_2 is
begin
-- TODO
end UB1BPPG_1_2;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_1_3 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_1_3;

architecture UB1BPPG_1_3 of UB1BPPG_1_3 is
begin
-- TODO
end UB1BPPG_1_3;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_1_4 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_1_4;

architecture UB1BPPG_1_4 of UB1BPPG_1_4 is
begin
-- TODO
end UB1BPPG_1_4;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_1_5 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_1_5;

architecture UB1BPPG_1_5 of UB1BPPG_1_5 is
begin
-- TODO
end UB1BPPG_1_5;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_1_6 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_1_6;

architecture UB1BPPG_1_6 of UB1BPPG_1_6 is
begin
-- TODO
end UB1BPPG_1_6;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_1_7 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_1_7;

architecture UB1BPPG_1_7 of UB1BPPG_1_7 is
begin
-- TODO
end UB1BPPG_1_7;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_2_0 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_2_0;

architecture UB1BPPG_2_0 of UB1BPPG_2_0 is
begin
-- TODO
end UB1BPPG_2_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_2_1 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_2_1;

architecture UB1BPPG_2_1 of UB1BPPG_2_1 is
begin
-- TODO
end UB1BPPG_2_1;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_2_2 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_2_2;

architecture UB1BPPG_2_2 of UB1BPPG_2_2 is
begin
-- TODO
end UB1BPPG_2_2;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_2_3 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_2_3;

architecture UB1BPPG_2_3 of UB1BPPG_2_3 is
begin
-- TODO
end UB1BPPG_2_3;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_2_4 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_2_4;

architecture UB1BPPG_2_4 of UB1BPPG_2_4 is
begin
-- TODO
end UB1BPPG_2_4;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_2_5 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_2_5;

architecture UB1BPPG_2_5 of UB1BPPG_2_5 is
begin
-- TODO
end UB1BPPG_2_5;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_2_6 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_2_6;

architecture UB1BPPG_2_6 of UB1BPPG_2_6 is
begin
-- TODO
end UB1BPPG_2_6;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_2_7 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_2_7;

architecture UB1BPPG_2_7 of UB1BPPG_2_7 is
begin
-- TODO
end UB1BPPG_2_7;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_3_0 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_3_0;

architecture UB1BPPG_3_0 of UB1BPPG_3_0 is
begin
-- TODO
end UB1BPPG_3_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_3_1 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_3_1;

architecture UB1BPPG_3_1 of UB1BPPG_3_1 is
begin
-- TODO
end UB1BPPG_3_1;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_3_2 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_3_2;

architecture UB1BPPG_3_2 of UB1BPPG_3_2 is
begin
-- TODO
end UB1BPPG_3_2;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_3_3 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_3_3;

architecture UB1BPPG_3_3 of UB1BPPG_3_3 is
begin
-- TODO
end UB1BPPG_3_3;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_3_4 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_3_4;

architecture UB1BPPG_3_4 of UB1BPPG_3_4 is
begin
-- TODO
end UB1BPPG_3_4;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_3_5 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_3_5;

architecture UB1BPPG_3_5 of UB1BPPG_3_5 is
begin
-- TODO
end UB1BPPG_3_5;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_3_6 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_3_6;

architecture UB1BPPG_3_6 of UB1BPPG_3_6 is
begin
-- TODO
end UB1BPPG_3_6;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_3_7 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_3_7;

architecture UB1BPPG_3_7 of UB1BPPG_3_7 is
begin
-- TODO
end UB1BPPG_3_7;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_4_0 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_4_0;

architecture UB1BPPG_4_0 of UB1BPPG_4_0 is
begin
-- TODO
end UB1BPPG_4_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_4_1 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_4_1;

architecture UB1BPPG_4_1 of UB1BPPG_4_1 is
begin
-- TODO
end UB1BPPG_4_1;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_4_2 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_4_2;

architecture UB1BPPG_4_2 of UB1BPPG_4_2 is
begin
-- TODO
end UB1BPPG_4_2;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_4_3 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_4_3;

architecture UB1BPPG_4_3 of UB1BPPG_4_3 is
begin
-- TODO
end UB1BPPG_4_3;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_4_4 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_4_4;

architecture UB1BPPG_4_4 of UB1BPPG_4_4 is
begin
-- TODO
end UB1BPPG_4_4;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_4_5 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_4_5;

architecture UB1BPPG_4_5 of UB1BPPG_4_5 is
begin
-- TODO
end UB1BPPG_4_5;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_4_6 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_4_6;

architecture UB1BPPG_4_6 of UB1BPPG_4_6 is
begin
-- TODO
end UB1BPPG_4_6;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_4_7 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_4_7;

architecture UB1BPPG_4_7 of UB1BPPG_4_7 is
begin
-- TODO
end UB1BPPG_4_7;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_5_0 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_5_0;

architecture UB1BPPG_5_0 of UB1BPPG_5_0 is
begin
-- TODO
end UB1BPPG_5_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_5_1 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_5_1;

architecture UB1BPPG_5_1 of UB1BPPG_5_1 is
begin
-- TODO
end UB1BPPG_5_1;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_5_2 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_5_2;

architecture UB1BPPG_5_2 of UB1BPPG_5_2 is
begin
-- TODO
end UB1BPPG_5_2;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_5_3 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_5_3;

architecture UB1BPPG_5_3 of UB1BPPG_5_3 is
begin
-- TODO
end UB1BPPG_5_3;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_5_4 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_5_4;

architecture UB1BPPG_5_4 of UB1BPPG_5_4 is
begin
-- TODO
end UB1BPPG_5_4;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_5_5 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_5_5;

architecture UB1BPPG_5_5 of UB1BPPG_5_5 is
begin
-- TODO
end UB1BPPG_5_5;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_5_6 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_5_6;

architecture UB1BPPG_5_6 of UB1BPPG_5_6 is
begin
-- TODO
end UB1BPPG_5_6;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_5_7 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_5_7;

architecture UB1BPPG_5_7 of UB1BPPG_5_7 is
begin
-- TODO
end UB1BPPG_5_7;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_6_0 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_6_0;

architecture UB1BPPG_6_0 of UB1BPPG_6_0 is
begin
-- TODO
end UB1BPPG_6_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_6_1 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_6_1;

architecture UB1BPPG_6_1 of UB1BPPG_6_1 is
begin
-- TODO
end UB1BPPG_6_1;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_6_2 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_6_2;

architecture UB1BPPG_6_2 of UB1BPPG_6_2 is
begin
-- TODO
end UB1BPPG_6_2;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_6_3 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_6_3;

architecture UB1BPPG_6_3 of UB1BPPG_6_3 is
begin
-- TODO
end UB1BPPG_6_3;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_6_4 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_6_4;

architecture UB1BPPG_6_4 of UB1BPPG_6_4 is
begin
-- TODO
end UB1BPPG_6_4;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_6_5 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_6_5;

architecture UB1BPPG_6_5 of UB1BPPG_6_5 is
begin
-- TODO
end UB1BPPG_6_5;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_6_6 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_6_6;

architecture UB1BPPG_6_6 of UB1BPPG_6_6 is
begin
-- TODO
end UB1BPPG_6_6;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_6_7 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_6_7;

architecture UB1BPPG_6_7 of UB1BPPG_6_7 is
begin
-- TODO
end UB1BPPG_6_7;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_7_0 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_7_0;

architecture UB1BPPG_7_0 of UB1BPPG_7_0 is
begin
-- TODO
end UB1BPPG_7_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_7_1 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_7_1;

architecture UB1BPPG_7_1 of UB1BPPG_7_1 is
begin
-- TODO
end UB1BPPG_7_1;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_7_2 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_7_2;

architecture UB1BPPG_7_2 of UB1BPPG_7_2 is
begin
-- TODO
end UB1BPPG_7_2;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_7_3 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_7_3;

architecture UB1BPPG_7_3 of UB1BPPG_7_3 is
begin
-- TODO
end UB1BPPG_7_3;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_7_4 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_7_4;

architecture UB1BPPG_7_4 of UB1BPPG_7_4 is
begin
-- TODO
end UB1BPPG_7_4;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_7_5 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_7_5;

architecture UB1BPPG_7_5 of UB1BPPG_7_5 is
begin
-- TODO
end UB1BPPG_7_5;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_7_6 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_7_6;

architecture UB1BPPG_7_6 of UB1BPPG_7_6 is
begin
-- TODO
end UB1BPPG_7_6;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1BPPG_7_7 is
  port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
end UB1BPPG_7_7;

architecture UB1BPPG_7_7 of UB1BPPG_7_7 is
begin
-- TODO
end UB1BPPG_7_7;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1DCON_0 is
  port(
      O : out std_logic;
      I : in std_logic);
end UB1DCON_0;

architecture UB1DCON_0 of UB1DCON_0 is
begin
-- TODO
end UB1DCON_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1DCON_1 is
  port(
      O : out std_logic;
      I : in std_logic);
end UB1DCON_1;

architecture UB1DCON_1 of UB1DCON_1 is
begin
-- TODO
end UB1DCON_1;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1DCON_10 is
  port(
      O : out std_logic;
      I : in std_logic);
end UB1DCON_10;

architecture UB1DCON_10 of UB1DCON_10 is
begin
-- TODO
end UB1DCON_10;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1DCON_11 is
  port(
      O : out std_logic;
      I : in std_logic);
end UB1DCON_11;

architecture UB1DCON_11 of UB1DCON_11 is
begin
-- TODO
end UB1DCON_11;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1DCON_12 is
  port(
      O : out std_logic;
      I : in std_logic);
end UB1DCON_12;

architecture UB1DCON_12 of UB1DCON_12 is
begin
-- TODO
end UB1DCON_12;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1DCON_13 is
  port(
      O : out std_logic;
      I : in std_logic);
end UB1DCON_13;

architecture UB1DCON_13 of UB1DCON_13 is
begin
-- TODO
end UB1DCON_13;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1DCON_14 is
  port(
      O : out std_logic;
      I : in std_logic);
end UB1DCON_14;

architecture UB1DCON_14 of UB1DCON_14 is
begin
-- TODO
end UB1DCON_14;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1DCON_2 is
  port(
      O : out std_logic;
      I : in std_logic);
end UB1DCON_2;

architecture UB1DCON_2 of UB1DCON_2 is
begin
-- TODO
end UB1DCON_2;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1DCON_3 is
  port(
      O : out std_logic;
      I : in std_logic);
end UB1DCON_3;

architecture UB1DCON_3 of UB1DCON_3 is
begin
-- TODO
end UB1DCON_3;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1DCON_4 is
  port(
      O : out std_logic;
      I : in std_logic);
end UB1DCON_4;

architecture UB1DCON_4 of UB1DCON_4 is
begin
-- TODO
end UB1DCON_4;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1DCON_5 is
  port(
      O : out std_logic;
      I : in std_logic);
end UB1DCON_5;

architecture UB1DCON_5 of UB1DCON_5 is
begin
-- TODO
end UB1DCON_5;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1DCON_6 is
  port(
      O : out std_logic;
      I : in std_logic);
end UB1DCON_6;

architecture UB1DCON_6 of UB1DCON_6 is
begin
-- TODO
end UB1DCON_6;

library IEEE;
use IEEE.std_logic_1164.all;
entity UB1DCON_9 is
  port(
      O : out std_logic;
      I : in std_logic);
end UB1DCON_9;

architecture UB1DCON_9 of UB1DCON_9 is
begin
-- TODO
end UB1DCON_9;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBARYACC_7_0_8_1_000 is
  port(
      S1 : out std_logic_vector(14 downto 7);
      S2 : out std_logic_vector(14 downto 0);
      PP0 : in std_logic_vector(7 downto 0);
      PP1 : in std_logic_vector(8 downto 1);
      PP2 : in std_logic_vector(9 downto 2);
      PP3 : in std_logic_vector(10 downto 3);
      PP4 : in std_logic_vector(11 downto 4);
      PP5 : in std_logic_vector(12 downto 5);
      PP6 : in std_logic_vector(13 downto 6);
      PP7 : in std_logic_vector(14 downto 7));
end UBARYACC_7_0_8_1_000;

architecture UBARYACC_7_0_8_1_000 of UBARYACC_7_0_8_1_000 is
  component CSA_7_0_8_1_9_2 
    port(
      C : out std_logic_vector(9 downto 2);
      S : out std_logic_vector(9 downto 0);
      X : in std_logic_vector(7 downto 0);
      Y : in std_logic_vector(8 downto 1);
      Z : in std_logic_vector(9 downto 2));
  end component;
  component CSA_9_0_9_2_10_3 
    port(
      C : out std_logic_vector(10 downto 3);
      S : out std_logic_vector(10 downto 0);
      X : in std_logic_vector(9 downto 0);
      Y : in std_logic_vector(9 downto 2);
      Z : in std_logic_vector(10 downto 3));
  end component;
  component CSA_10_0_10_3_11_000 
    port(
      C : out std_logic_vector(11 downto 4);
      S : out std_logic_vector(11 downto 0);
      X : in std_logic_vector(10 downto 0);
      Y : in std_logic_vector(10 downto 3);
      Z : in std_logic_vector(11 downto 4));
  end component;
  component CSA_11_0_11_4_12_000 
    port(
      C : out std_logic_vector(12 downto 5);
      S : out std_logic_vector(12 downto 0);
      X : in std_logic_vector(11 downto 0);
      Y : in std_logic_vector(11 downto 4);
      Z : in std_logic_vector(12 downto 5));
  end component;
  component CSA_12_0_12_5_13_000 
    port(
      C : out std_logic_vector(13 downto 6);
      S : out std_logic_vector(13 downto 0);
      X : in std_logic_vector(12 downto 0);
      Y : in std_logic_vector(12 downto 5);
      Z : in std_logic_vector(13 downto 6));
  end component;
  component CSA_13_0_13_6_14_000 
    port(
      C : out std_logic_vector(14 downto 7);
      S : out std_logic_vector(14 downto 0);
      X : in std_logic_vector(13 downto 0);
      Y : in std_logic_vector(13 downto 6);
      Z : in std_logic_vector(14 downto 7));
  end component;
  signal IC0 : std_logic_vector(9 downto 2);
  signal IC1 : std_logic_vector(10 downto 3);
  signal IC2 : std_logic_vector(11 downto 4);
  signal IC3 : std_logic_vector(12 downto 5);
  signal IC4 : std_logic_vector(13 downto 6);
  signal IS0 : std_logic_vector(9 downto 0);
  signal IS1 : std_logic_vector(10 downto 0);
  signal IS2 : std_logic_vector(11 downto 0);
  signal IS3 : std_logic_vector(12 downto 0);
  signal IS4 : std_logic_vector(13 downto 0);
begin
  U0: CSA_7_0_8_1_9_2 port map (IC0, IS0, PP0, PP1, PP2);
  U1: CSA_9_0_9_2_10_3 port map (IC1, IS1, IS0, IC0, PP3);
  U2: CSA_10_0_10_3_11_000 port map (IC2, IS2, IS1, IC1, PP4);
  U3: CSA_11_0_11_4_12_000 port map (IC3, IS3, IS2, IC2, PP5);
  U4: CSA_12_0_12_5_13_000 port map (IC4, IS4, IS3, IC3, PP6);
  U5: CSA_13_0_13_6_14_000 port map (S1, S2, IS4, IC4, PP7);
end UBARYACC_7_0_8_1_000;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBCON_1_0 is
  port(
      O : out std_logic_vector(1 downto 0);
      I : in std_logic_vector(1 downto 0));
end UBCON_1_0;

architecture UBCON_1_0 of UBCON_1_0 is
  component UB1DCON_0 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_1 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
begin
  U0: UB1DCON_0 port map (O(0), I(0));
  U1: UB1DCON_1 port map (O(1), I(1));
end UBCON_1_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBCON_2_0 is
  port(
      O : out std_logic_vector(2 downto 0);
      I : in std_logic_vector(2 downto 0));
end UBCON_2_0;

architecture UBCON_2_0 of UBCON_2_0 is
  component UB1DCON_0 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_1 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_2 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
begin
  U0: UB1DCON_0 port map (O(0), I(0));
  U1: UB1DCON_1 port map (O(1), I(1));
  U2: UB1DCON_2 port map (O(2), I(2));
end UBCON_2_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBCON_3_0 is
  port(
      O : out std_logic_vector(3 downto 0);
      I : in std_logic_vector(3 downto 0));
end UBCON_3_0;

architecture UBCON_3_0 of UBCON_3_0 is
  component UB1DCON_0 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_1 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_2 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_3 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
begin
  U0: UB1DCON_0 port map (O(0), I(0));
  U1: UB1DCON_1 port map (O(1), I(1));
  U2: UB1DCON_2 port map (O(2), I(2));
  U3: UB1DCON_3 port map (O(3), I(3));
end UBCON_3_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBCON_4_0 is
  port(
      O : out std_logic_vector(4 downto 0);
      I : in std_logic_vector(4 downto 0));
end UBCON_4_0;

architecture UBCON_4_0 of UBCON_4_0 is
  component UB1DCON_0 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_1 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_2 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_3 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_4 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
begin
  U0: UB1DCON_0 port map (O(0), I(0));
  U1: UB1DCON_1 port map (O(1), I(1));
  U2: UB1DCON_2 port map (O(2), I(2));
  U3: UB1DCON_3 port map (O(3), I(3));
  U4: UB1DCON_4 port map (O(4), I(4));
end UBCON_4_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBCON_5_0 is
  port(
      O : out std_logic_vector(5 downto 0);
      I : in std_logic_vector(5 downto 0));
end UBCON_5_0;

architecture UBCON_5_0 of UBCON_5_0 is
  component UB1DCON_0 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_1 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_2 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_3 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_4 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_5 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
begin
  U0: UB1DCON_0 port map (O(0), I(0));
  U1: UB1DCON_1 port map (O(1), I(1));
  U2: UB1DCON_2 port map (O(2), I(2));
  U3: UB1DCON_3 port map (O(3), I(3));
  U4: UB1DCON_4 port map (O(4), I(4));
  U5: UB1DCON_5 port map (O(5), I(5));
end UBCON_5_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBCON_6_0 is
  port(
      O : out std_logic_vector(6 downto 0);
      I : in std_logic_vector(6 downto 0));
end UBCON_6_0;

architecture UBCON_6_0 of UBCON_6_0 is
  component UB1DCON_0 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_1 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_2 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_3 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_4 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_5 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
  component UB1DCON_6 
    port(
      O : out std_logic;
      I : in std_logic);
  end component;
begin
  U0: UB1DCON_0 port map (O(0), I(0));
  U1: UB1DCON_1 port map (O(1), I(1));
  U2: UB1DCON_2 port map (O(2), I(2));
  U3: UB1DCON_3 port map (O(3), I(3));
  U4: UB1DCON_4 port map (O(4), I(4));
  U5: UB1DCON_5 port map (O(5), I(5));
  U6: UB1DCON_6 port map (O(6), I(6));
end UBCON_6_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBFA_10 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
end UBFA_10;

architecture UBFA_10 of UBFA_10 is
begin
-- TODO
end UBFA_10;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBFA_11 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
end UBFA_11;

architecture UBFA_11 of UBFA_11 is
begin
-- TODO
end UBFA_11;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBFA_12 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
end UBFA_12;

architecture UBFA_12 of UBFA_12 is
begin
-- TODO
end UBFA_12;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBFA_13 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
end UBFA_13;

architecture UBFA_13 of UBFA_13 is
begin
-- TODO
end UBFA_13;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBFA_2 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
end UBFA_2;

architecture UBFA_2 of UBFA_2 is
begin
-- TODO
end UBFA_2;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBFA_3 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
end UBFA_3;

architecture UBFA_3 of UBFA_3 is
begin
-- TODO
end UBFA_3;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBFA_4 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
end UBFA_4;

architecture UBFA_4 of UBFA_4 is
begin
-- TODO
end UBFA_4;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBFA_5 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
end UBFA_5;

architecture UBFA_5 of UBFA_5 is
begin
-- TODO
end UBFA_5;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBFA_6 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
end UBFA_6;

architecture UBFA_6 of UBFA_6 is
begin
-- TODO
end UBFA_6;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBFA_7 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
end UBFA_7;

architecture UBFA_7 of UBFA_7 is
begin
-- TODO
end UBFA_7;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBFA_8 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
end UBFA_8;

architecture UBFA_8 of UBFA_8 is
begin
-- TODO
end UBFA_8;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBFA_9 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic;
      Z : in std_logic);
end UBFA_9;

architecture UBFA_9 of UBFA_9 is
begin
-- TODO
end UBFA_9;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBHA_1 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic);
end UBHA_1;

architecture UBHA_1 of UBHA_1 is
begin
-- TODO
end UBHA_1;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBHA_2 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic);
end UBHA_2;

architecture UBHA_2 of UBHA_2 is
begin
-- TODO
end UBHA_2;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBHA_3 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic);
end UBHA_3;

architecture UBHA_3 of UBHA_3 is
begin
-- TODO
end UBHA_3;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBHA_4 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic);
end UBHA_4;

architecture UBHA_4 of UBHA_4 is
begin
-- TODO
end UBHA_4;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBHA_5 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic);
end UBHA_5;

architecture UBHA_5 of UBHA_5 is
begin
-- TODO
end UBHA_5;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBHA_6 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic);
end UBHA_6;

architecture UBHA_6 of UBHA_6 is
begin
-- TODO
end UBHA_6;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBHA_8 is
  port(
      C : out std_logic;
      S : out std_logic;
      X : in std_logic;
      Y : in std_logic);
end UBHA_8;

architecture UBHA_8 of UBHA_8 is
begin
-- TODO
end UBHA_8;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBHCA_14_7_14_0 is
  port(
      S : out std_logic_vector(15 downto 0);
      X : in std_logic_vector(14 downto 7);
      Y : in std_logic_vector(14 downto 0));
end UBHCA_14_7_14_0;

architecture UBHCA_14_7_14_0 of UBHCA_14_7_14_0 is
  component UBPureHCA_14_7 
    port(
      S : out std_logic_vector(15 downto 7);
      X : in std_logic_vector(14 downto 7);
      Y : in std_logic_vector(14 downto 7));
  end component;
  component UBCON_6_0 
    port(
      O : out std_logic_vector(6 downto 0);
      I : in std_logic_vector(6 downto 0));
  end component;
begin
  U0: UBPureHCA_14_7 port map (S(15 downto 7), X(14 downto 7), Y(14 downto 7));
  U1: UBCON_6_0 port map (S(6 downto 0), Y(6 downto 0));
end UBHCA_14_7_14_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBPPG_7_0_7_0 is
  port(
      PP0 : out std_logic_vector(7 downto 0);
      PP1 : out std_logic_vector(8 downto 1);
      PP2 : out std_logic_vector(9 downto 2);
      PP3 : out std_logic_vector(10 downto 3);
      PP4 : out std_logic_vector(11 downto 4);
      PP5 : out std_logic_vector(12 downto 5);
      PP6 : out std_logic_vector(13 downto 6);
      PP7 : out std_logic_vector(14 downto 7);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic_vector(7 downto 0));
end UBPPG_7_0_7_0;

architecture UBPPG_7_0_7_0 of UBPPG_7_0_7_0 is
  component UBVPPG_7_0_0 
    port(
      O : out std_logic_vector(7 downto 0);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
  end component;
  component UBVPPG_7_0_1 
    port(
      O : out std_logic_vector(8 downto 1);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
  end component;
  component UBVPPG_7_0_2 
    port(
      O : out std_logic_vector(9 downto 2);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
  end component;
  component UBVPPG_7_0_3 
    port(
      O : out std_logic_vector(10 downto 3);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
  end component;
  component UBVPPG_7_0_4 
    port(
      O : out std_logic_vector(11 downto 4);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
  end component;
  component UBVPPG_7_0_5 
    port(
      O : out std_logic_vector(12 downto 5);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
  end component;
  component UBVPPG_7_0_6 
    port(
      O : out std_logic_vector(13 downto 6);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
  end component;
  component UBVPPG_7_0_7 
    port(
      O : out std_logic_vector(14 downto 7);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
  end component;
begin
  U0: UBVPPG_7_0_0 port map (PP0, IN1, IN2(0));
  U1: UBVPPG_7_0_1 port map (PP1, IN1, IN2(1));
  U2: UBVPPG_7_0_2 port map (PP2, IN1, IN2(2));
  U3: UBVPPG_7_0_3 port map (PP3, IN1, IN2(3));
  U4: UBVPPG_7_0_4 port map (PP4, IN1, IN2(4));
  U5: UBVPPG_7_0_5 port map (PP5, IN1, IN2(5));
  U6: UBVPPG_7_0_6 port map (PP6, IN1, IN2(6));
  U7: UBVPPG_7_0_7 port map (PP7, IN1, IN2(7));
end UBPPG_7_0_7_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBPriHCA_14_7 is
  port(
      S : out std_logic_vector(15 downto 7);
      X : in std_logic_vector(14 downto 7);
      Y : in std_logic_vector(14 downto 7);
      Cin : in std_logic);
end UBPriHCA_14_7;

architecture UBPriHCA_14_7 of UBPriHCA_14_7 is
begin
-- TODO
end UBPriHCA_14_7;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBPureHCA_14_7 is
  port(
      S : out std_logic_vector(15 downto 7);
      X : in std_logic_vector(14 downto 7);
      Y : in std_logic_vector(14 downto 7));
end UBPureHCA_14_7;

architecture UBPureHCA_14_7 of UBPureHCA_14_7 is
  component UBPriHCA_14_7 
    port(
      S : out std_logic_vector(15 downto 7);
      X : in std_logic_vector(14 downto 7);
      Y : in std_logic_vector(14 downto 7);
      Cin : in std_logic);
  end component;
  component UBZero_7_7 
    port(
      O : out std_logic);
  end component;
  signal C : std_logic;
begin
  U0: UBPriHCA_14_7 port map (S, X, Y, C);
  U1: UBZero_7_7 port map (C);
end UBPureHCA_14_7;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBVPPG_7_0_0 is
  port(
      O : out std_logic_vector(7 downto 0);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
end UBVPPG_7_0_0;

architecture UBVPPG_7_0_0 of UBVPPG_7_0_0 is
  component UB1BPPG_0_0 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_1_0 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_2_0 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_3_0 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_4_0 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_5_0 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_6_0 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_7_0 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
begin
  U0: UB1BPPG_0_0 port map (O(0), IN1(0), IN2);
  U1: UB1BPPG_1_0 port map (O(1), IN1(1), IN2);
  U2: UB1BPPG_2_0 port map (O(2), IN1(2), IN2);
  U3: UB1BPPG_3_0 port map (O(3), IN1(3), IN2);
  U4: UB1BPPG_4_0 port map (O(4), IN1(4), IN2);
  U5: UB1BPPG_5_0 port map (O(5), IN1(5), IN2);
  U6: UB1BPPG_6_0 port map (O(6), IN1(6), IN2);
  U7: UB1BPPG_7_0 port map (O(7), IN1(7), IN2);
end UBVPPG_7_0_0;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBVPPG_7_0_1 is
  port(
      O : out std_logic_vector(8 downto 1);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
end UBVPPG_7_0_1;

architecture UBVPPG_7_0_1 of UBVPPG_7_0_1 is
  component UB1BPPG_0_1 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_1_1 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_2_1 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_3_1 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_4_1 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_5_1 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_6_1 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_7_1 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
begin
  U0: UB1BPPG_0_1 port map (O(1), IN1(0), IN2);
  U1: UB1BPPG_1_1 port map (O(2), IN1(1), IN2);
  U2: UB1BPPG_2_1 port map (O(3), IN1(2), IN2);
  U3: UB1BPPG_3_1 port map (O(4), IN1(3), IN2);
  U4: UB1BPPG_4_1 port map (O(5), IN1(4), IN2);
  U5: UB1BPPG_5_1 port map (O(6), IN1(5), IN2);
  U6: UB1BPPG_6_1 port map (O(7), IN1(6), IN2);
  U7: UB1BPPG_7_1 port map (O(8), IN1(7), IN2);
end UBVPPG_7_0_1;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBVPPG_7_0_2 is
  port(
      O : out std_logic_vector(9 downto 2);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
end UBVPPG_7_0_2;

architecture UBVPPG_7_0_2 of UBVPPG_7_0_2 is
  component UB1BPPG_0_2 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_1_2 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_2_2 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_3_2 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_4_2 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_5_2 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_6_2 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_7_2 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
begin
  U0: UB1BPPG_0_2 port map (O(2), IN1(0), IN2);
  U1: UB1BPPG_1_2 port map (O(3), IN1(1), IN2);
  U2: UB1BPPG_2_2 port map (O(4), IN1(2), IN2);
  U3: UB1BPPG_3_2 port map (O(5), IN1(3), IN2);
  U4: UB1BPPG_4_2 port map (O(6), IN1(4), IN2);
  U5: UB1BPPG_5_2 port map (O(7), IN1(5), IN2);
  U6: UB1BPPG_6_2 port map (O(8), IN1(6), IN2);
  U7: UB1BPPG_7_2 port map (O(9), IN1(7), IN2);
end UBVPPG_7_0_2;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBVPPG_7_0_3 is
  port(
      O : out std_logic_vector(10 downto 3);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
end UBVPPG_7_0_3;

architecture UBVPPG_7_0_3 of UBVPPG_7_0_3 is
  component UB1BPPG_0_3 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_1_3 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_2_3 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_3_3 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_4_3 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_5_3 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_6_3 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_7_3 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
begin
  U0: UB1BPPG_0_3 port map (O(3), IN1(0), IN2);
  U1: UB1BPPG_1_3 port map (O(4), IN1(1), IN2);
  U2: UB1BPPG_2_3 port map (O(5), IN1(2), IN2);
  U3: UB1BPPG_3_3 port map (O(6), IN1(3), IN2);
  U4: UB1BPPG_4_3 port map (O(7), IN1(4), IN2);
  U5: UB1BPPG_5_3 port map (O(8), IN1(5), IN2);
  U6: UB1BPPG_6_3 port map (O(9), IN1(6), IN2);
  U7: UB1BPPG_7_3 port map (O(10), IN1(7), IN2);
end UBVPPG_7_0_3;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBVPPG_7_0_4 is
  port(
      O : out std_logic_vector(11 downto 4);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
end UBVPPG_7_0_4;

architecture UBVPPG_7_0_4 of UBVPPG_7_0_4 is
  component UB1BPPG_0_4 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_1_4 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_2_4 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_3_4 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_4_4 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_5_4 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_6_4 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_7_4 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
begin
  U0: UB1BPPG_0_4 port map (O(4), IN1(0), IN2);
  U1: UB1BPPG_1_4 port map (O(5), IN1(1), IN2);
  U2: UB1BPPG_2_4 port map (O(6), IN1(2), IN2);
  U3: UB1BPPG_3_4 port map (O(7), IN1(3), IN2);
  U4: UB1BPPG_4_4 port map (O(8), IN1(4), IN2);
  U5: UB1BPPG_5_4 port map (O(9), IN1(5), IN2);
  U6: UB1BPPG_6_4 port map (O(10), IN1(6), IN2);
  U7: UB1BPPG_7_4 port map (O(11), IN1(7), IN2);
end UBVPPG_7_0_4;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBVPPG_7_0_5 is
  port(
      O : out std_logic_vector(12 downto 5);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
end UBVPPG_7_0_5;

architecture UBVPPG_7_0_5 of UBVPPG_7_0_5 is
  component UB1BPPG_0_5 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_1_5 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_2_5 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_3_5 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_4_5 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_5_5 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_6_5 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_7_5 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
begin
  U0: UB1BPPG_0_5 port map (O(5), IN1(0), IN2);
  U1: UB1BPPG_1_5 port map (O(6), IN1(1), IN2);
  U2: UB1BPPG_2_5 port map (O(7), IN1(2), IN2);
  U3: UB1BPPG_3_5 port map (O(8), IN1(3), IN2);
  U4: UB1BPPG_4_5 port map (O(9), IN1(4), IN2);
  U5: UB1BPPG_5_5 port map (O(10), IN1(5), IN2);
  U6: UB1BPPG_6_5 port map (O(11), IN1(6), IN2);
  U7: UB1BPPG_7_5 port map (O(12), IN1(7), IN2);
end UBVPPG_7_0_5;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBVPPG_7_0_6 is
  port(
      O : out std_logic_vector(13 downto 6);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
end UBVPPG_7_0_6;

architecture UBVPPG_7_0_6 of UBVPPG_7_0_6 is
  component UB1BPPG_0_6 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_1_6 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_2_6 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_3_6 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_4_6 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_5_6 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_6_6 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_7_6 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
begin
  U0: UB1BPPG_0_6 port map (O(6), IN1(0), IN2);
  U1: UB1BPPG_1_6 port map (O(7), IN1(1), IN2);
  U2: UB1BPPG_2_6 port map (O(8), IN1(2), IN2);
  U3: UB1BPPG_3_6 port map (O(9), IN1(3), IN2);
  U4: UB1BPPG_4_6 port map (O(10), IN1(4), IN2);
  U5: UB1BPPG_5_6 port map (O(11), IN1(5), IN2);
  U6: UB1BPPG_6_6 port map (O(12), IN1(6), IN2);
  U7: UB1BPPG_7_6 port map (O(13), IN1(7), IN2);
end UBVPPG_7_0_6;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBVPPG_7_0_7 is
  port(
      O : out std_logic_vector(14 downto 7);
      IN1 : in std_logic_vector(7 downto 0);
      IN2 : in std_logic);
end UBVPPG_7_0_7;

architecture UBVPPG_7_0_7 of UBVPPG_7_0_7 is
  component UB1BPPG_0_7 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_1_7 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_2_7 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_3_7 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_4_7 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_5_7 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_6_7 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
  component UB1BPPG_7_7 
    port(
      O : out std_logic;
      IN1 : in std_logic;
      IN2 : in std_logic);
  end component;
begin
  U0: UB1BPPG_0_7 port map (O(7), IN1(0), IN2);
  U1: UB1BPPG_1_7 port map (O(8), IN1(1), IN2);
  U2: UB1BPPG_2_7 port map (O(9), IN1(2), IN2);
  U3: UB1BPPG_3_7 port map (O(10), IN1(3), IN2);
  U4: UB1BPPG_4_7 port map (O(11), IN1(4), IN2);
  U5: UB1BPPG_5_7 port map (O(12), IN1(5), IN2);
  U6: UB1BPPG_6_7 port map (O(13), IN1(6), IN2);
  U7: UB1BPPG_7_7 port map (O(14), IN1(7), IN2);
end UBVPPG_7_0_7;

library IEEE;
use IEEE.std_logic_1164.all;
entity UBZero_7_7 is
  port(
      O : out std_logic);
end UBZero_7_7;

architecture UBZero_7_7 of UBZero_7_7 is
begin
-- TODO
end UBZero_7_7;

