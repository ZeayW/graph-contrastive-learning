/*----------------------------------------------------------------------------
  Copyright (c) 2021 Homma laboratory. All rights reserved.

  Top module: Multiplier_13_0_1000

  Number system: Unsigned binary
  Multiplicand length: 14
  Multiplier length: 14
  Partial product generation: Simple PPG
  Partial product accumulation: Overturned-stairs tree
  Final stage addition: Carry select adder
----------------------------------------------------------------------------*/

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_1(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_2(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_12(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_13(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_14(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_14(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_15(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_16(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_17(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_7(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_17(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_18(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_19(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_20(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_21(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_6(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_19(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_21(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_5(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_18(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_10(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_20(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_21(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_22(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_23(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_24(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_11(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_23(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_24(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB1DCON_25(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_9(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_22(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_24(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_25(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_8(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_23(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_12(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_25(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_26(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBZero_27_27(O);
  output [27:27] O;
  assign O[27] = 0;
endmodule

module UBOne_6(O);
  output O;
  assign O = 1;
endmodule

module UBZero_6_6(O);
  output [6:6] O;
  assign O[6] = 0;
endmodule

module UBCSlB_6_6(Co, S, X, Y, Ci);
  output Co;
  output [6:6] S;
  input Ci;
  input [6:6] X;
  input [6:6] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [6:6] S_0;
  wire [6:6] S_1;
  assign S[6] = ( S_0[6] & ( ~ Ci ) ) | ( S_1[6] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_6 U0 (Ci_1);
  UBZero_6_6 U1 (Ci_0);
  UBRCB_6_6 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_6_6 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_7(O);
  output O;
  assign O = 1;
endmodule

module UBZero_7_7(O);
  output [7:7] O;
  assign O[7] = 0;
endmodule

module UBCSlB_8_7(Co, S, X, Y, Ci);
  output Co;
  output [8:7] S;
  input Ci;
  input [8:7] X;
  input [8:7] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [8:7] S_0;
  wire [8:7] S_1;
  assign S[7] = ( S_0[7] & ( ~ Ci ) ) | ( S_1[7] & Ci );
  assign S[8] = ( S_0[8] & ( ~ Ci ) ) | ( S_1[8] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_7 U0 (Ci_1);
  UBZero_7_7 U1 (Ci_0);
  UBRCB_8_7 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_8_7 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_9(O);
  output O;
  assign O = 1;
endmodule

module UBZero_9_9(O);
  output [9:9] O;
  assign O[9] = 0;
endmodule

module UBCSlB_11_9(Co, S, X, Y, Ci);
  output Co;
  output [11:9] S;
  input Ci;
  input [11:9] X;
  input [11:9] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [11:9] S_0;
  wire [11:9] S_1;
  assign S[9] = ( S_0[9] & ( ~ Ci ) ) | ( S_1[9] & Ci );
  assign S[10] = ( S_0[10] & ( ~ Ci ) ) | ( S_1[10] & Ci );
  assign S[11] = ( S_0[11] & ( ~ Ci ) ) | ( S_1[11] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_9 U0 (Ci_1);
  UBZero_9_9 U1 (Ci_0);
  UBRCB_11_9 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_11_9 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_12(O);
  output O;
  assign O = 1;
endmodule

module UBZero_12_12(O);
  output [12:12] O;
  assign O[12] = 0;
endmodule

module UBCSlB_15_12(Co, S, X, Y, Ci);
  output Co;
  output [15:12] S;
  input Ci;
  input [15:12] X;
  input [15:12] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [15:12] S_0;
  wire [15:12] S_1;
  assign S[12] = ( S_0[12] & ( ~ Ci ) ) | ( S_1[12] & Ci );
  assign S[13] = ( S_0[13] & ( ~ Ci ) ) | ( S_1[13] & Ci );
  assign S[14] = ( S_0[14] & ( ~ Ci ) ) | ( S_1[14] & Ci );
  assign S[15] = ( S_0[15] & ( ~ Ci ) ) | ( S_1[15] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_12 U0 (Ci_1);
  UBZero_12_12 U1 (Ci_0);
  UBRCB_15_12 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_15_12 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_16(O);
  output O;
  assign O = 1;
endmodule

module UBZero_16_16(O);
  output [16:16] O;
  assign O[16] = 0;
endmodule

module UBCSlB_20_16(Co, S, X, Y, Ci);
  output Co;
  output [20:16] S;
  input Ci;
  input [20:16] X;
  input [20:16] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [20:16] S_0;
  wire [20:16] S_1;
  assign S[16] = ( S_0[16] & ( ~ Ci ) ) | ( S_1[16] & Ci );
  assign S[17] = ( S_0[17] & ( ~ Ci ) ) | ( S_1[17] & Ci );
  assign S[18] = ( S_0[18] & ( ~ Ci ) ) | ( S_1[18] & Ci );
  assign S[19] = ( S_0[19] & ( ~ Ci ) ) | ( S_1[19] & Ci );
  assign S[20] = ( S_0[20] & ( ~ Ci ) ) | ( S_1[20] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_16 U0 (Ci_1);
  UBZero_16_16 U1 (Ci_0);
  UBRCB_20_16 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_20_16 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_21(O);
  output O;
  assign O = 1;
endmodule

module UBZero_21_21(O);
  output [21:21] O;
  assign O[21] = 0;
endmodule

module UBCSlB_26_21(Co, S, X, Y, Ci);
  output Co;
  output [26:21] S;
  input Ci;
  input [26:21] X;
  input [26:21] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [26:21] S_0;
  wire [26:21] S_1;
  assign S[21] = ( S_0[21] & ( ~ Ci ) ) | ( S_1[21] & Ci );
  assign S[22] = ( S_0[22] & ( ~ Ci ) ) | ( S_1[22] & Ci );
  assign S[23] = ( S_0[23] & ( ~ Ci ) ) | ( S_1[23] & Ci );
  assign S[24] = ( S_0[24] & ( ~ Ci ) ) | ( S_1[24] & Ci );
  assign S[25] = ( S_0[25] & ( ~ Ci ) ) | ( S_1[25] & Ci );
  assign S[26] = ( S_0[26] & ( ~ Ci ) ) | ( S_1[26] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_21 U0 (Ci_1);
  UBZero_21_21 U1 (Ci_0);
  UBRCB_26_21 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_26_21 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBOne_27(O);
  output O;
  assign O = 1;
endmodule

module UBFA_27(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBCSlB_27_27(Co, S, X, Y, Ci);
  output Co;
  output [27:27] S;
  input Ci;
  input [27:27] X;
  input [27:27] Y;
  wire Ci_0;
  wire Ci_1;
  wire Co_0;
  wire Co_1;
  wire [27:27] S_0;
  wire [27:27] S_1;
  assign S[27] = ( S_0[27] & ( ~ Ci ) ) | ( S_1[27] & Ci );
  assign Co = ( Co_0 & ( ~ Ci ) ) | ( Co_1 & Ci );
  UBOne_27 U0 (Ci_1);
  UBZero_27_27 U1 (Ci_0);
  UBRCB_27_27 U2 (Co_0, S_0, X, Y, Ci_0);
  UBRCB_27_27 U3 (Co_1, S_1, X, Y, Ci_1);
endmodule

module UBPriCSlA_27_5(S, X, Y, Cin);
  output [28:5] S;
  input Cin;
  input [27:5] X;
  input [27:5] Y;
  wire C0;
  wire C1;
  wire C2;
  wire C3;
  wire C4;
  wire C5;
  wire C6;
  UBRCB_5_5 U0 (C0, S[5], X[5], Y[5], Cin);
  UBCSlB_6_6 U1 (C1, S[6], X[6], Y[6], C0);
  UBCSlB_8_7 U2 (C2, S[8:7], X[8:7], Y[8:7], C1);
  UBCSlB_11_9 U3 (C3, S[11:9], X[11:9], Y[11:9], C2);
  UBCSlB_15_12 U4 (C4, S[15:12], X[15:12], Y[15:12], C3);
  UBCSlB_20_16 U5 (C5, S[20:16], X[20:16], Y[20:16], C4);
  UBCSlB_26_21 U6 (C6, S[26:21], X[26:21], Y[26:21], C5);
  UBCSlB_27_27 U7 (S[28], S[27], X[27], Y[27], C6);
endmodule

module UBZero_5_5(O);
  output [5:5] O;
  assign O[5] = 0;
endmodule

module Multiplier_13_0_1000(P, IN1, IN2);
  output [27:0] P;
  input [13:0] IN1;
  input [13:0] IN2;
  wire [28:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  assign P[12] = W[12];
  assign P[13] = W[13];
  assign P[14] = W[14];
  assign P[15] = W[15];
  assign P[16] = W[16];
  assign P[17] = W[17];
  assign P[18] = W[18];
  assign P[19] = W[19];
  assign P[20] = W[20];
  assign P[21] = W[21];
  assign P[22] = W[22];
  assign P[23] = W[23];
  assign P[24] = W[24];
  assign P[25] = W[25];
  assign P[26] = W[26];
  assign P[27] = W[27];
  MultUB_STD_OS_CSe000 U0 (W, IN1, IN2);
endmodule

module CSA_13_0_14_1_15_000 (C, S, X, Y, Z);
  output [15:2] C;
  output [15:0] S;
  input [13:0] X;
  input [14:1] Y;
  input [15:2] Z;
  UB1DCON_0 U0 (S[0], X[0]);
  UBHA_1 U1 (C[2], S[1], Y[1], X[1]);
  PureCSA_13_2 U2 (C[14:3], S[13:2], Z[13:2], Y[13:2], X[13:2]);
  UBHA_14 U3 (C[15], S[14], Z[14], Y[14]);
  UB1DCON_15 U4 (S[15], Z[15]);
endmodule

module CSA_15_2_15_0_18_000 (C, S, X, Y, Z);
  output [16:3] C;
  output [18:0] S;
  input [15:2] X;
  input [15:0] Y;
  input [18:5] Z;
  UBCON_1_0 U0 (S[1:0], Y[1:0]);
  PureCSHA_4_2 U1 (C[5:3], S[4:2], X[4:2], Y[4:2]);
  PureCSA_15_5 U2 (C[16:6], S[15:5], Z[15:5], X[15:5], Y[15:5]);
  UBCON_18_16 U3 (S[18:16], Z[18:16]);
endmodule

module CSA_16_3_17_4_18_000 (C, S, X, Y, Z);
  output [18:5] C;
  output [18:3] S;
  input [16:3] X;
  input [17:4] Y;
  input [18:5] Z;
  UB1DCON_3 U0 (S[3], X[3]);
  UBHA_4 U1 (C[5], S[4], Y[4], X[4]);
  PureCSA_16_5 U2 (C[17:6], S[16:5], Z[16:5], Y[16:5], X[16:5]);
  UBHA_17 U3 (C[18], S[17], Z[17], Y[17]);
  UB1DCON_18 U4 (S[18], Z[18]);
endmodule

module CSA_16_3_18_0_22_000 (C, S, X, Y, Z);
  output [19:4] C;
  output [22:0] S;
  input [16:3] X;
  input [18:0] Y;
  input [22:7] Z;
  UBCON_2_0 U0 (S[2:0], Y[2:0]);
  PureCSHA_6_3 U1 (C[7:4], S[6:3], X[6:3], Y[6:3]);
  PureCSA_16_7 U2 (C[17:8], S[16:7], Z[16:7], X[16:7], Y[16:7]);
  PureCSHA_18_17 U3 (C[19:18], S[18:17], Z[18:17], Y[18:17]);
  UBCON_22_19 U4 (S[22:19], Z[22:19]);
endmodule

module CSA_18_3_21_8_21_000 (C, S, X, Y, Z);
  output [22:7] C;
  output [21:3] S;
  input [18:3] X;
  input [21:8] Y;
  input [21:6] Z;
  UBCON_5_3 U0 (S[5:3], X[5:3]);
  PureCSHA_7_6 U1 (C[8:7], S[7:6], Z[7:6], X[7:6]);
  PureCSA_18_8 U2 (C[19:9], S[18:8], Y[18:8], Z[18:8], X[18:8]);
  PureCSHA_21_19 U3 (C[22:20], S[21:19], Z[21:19], Y[21:19]);
endmodule

module CSA_19_4_22_0_26_000 (C, S, X, Y, Z);
  output [23:5] C;
  output [26:0] S;
  input [19:4] X;
  input [22:0] Y;
  input [26:10] Z;
  UBCON_3_0 U0 (S[3:0], Y[3:0]);
  PureCSHA_9_4 U1 (C[10:5], S[9:4], X[9:4], Y[9:4]);
  PureCSA_19_10 U2 (C[20:11], S[19:10], Z[19:10], X[19:10], Y[19:10]);
  PureCSHA_22_20 U3 (C[23:21], S[22:20], Z[22:20], Y[22:20]);
  UBCON_26_23 U4 (S[26:23], Z[26:23]);
endmodule

module CSA_19_6_20_7_21_000 (C, S, X, Y, Z);
  output [21:8] C;
  output [21:6] S;
  input [19:6] X;
  input [20:7] Y;
  input [21:8] Z;
  UB1DCON_6 U0 (S[6], X[6]);
  UBHA_7 U1 (C[8], S[7], Y[7], X[7]);
  PureCSA_19_8 U2 (C[20:9], S[19:8], Z[19:8], Y[19:8], X[19:8]);
  UBHA_20 U3 (C[21], S[20], Z[20], Y[20]);
  UB1DCON_21 U4 (S[21], Z[21]);
endmodule

module CSA_21_3_25_12_25000 (C, S, X, Y, Z);
  output [26:10] C;
  output [25:3] S;
  input [21:3] X;
  input [25:12] Y;
  input [25:9] Z;
  UBCON_8_3 U0 (S[8:3], X[8:3]);
  PureCSHA_11_9 U1 (C[12:10], S[11:9], Z[11:9], X[11:9]);
  PureCSA_21_12 U2 (C[22:13], S[21:12], Y[21:12], Z[21:12], X[21:12]);
  PureCSHA_25_22 U3 (C[26:23], S[25:22], Z[25:22], Y[25:22]);
endmodule

module CSA_22_9_23_10_24000 (C, S, X, Y, Z);
  output [24:11] C;
  output [24:9] S;
  input [22:9] X;
  input [23:10] Y;
  input [24:11] Z;
  UB1DCON_9 U0 (S[9], X[9]);
  UBHA_10 U1 (C[11], S[10], Y[10], X[10]);
  PureCSA_22_11 U2 (C[23:12], S[22:11], Z[22:11], Y[22:11], X[22:11]);
  UBHA_23 U3 (C[24], S[23], Z[23], Y[23]);
  UB1DCON_24 U4 (S[24], Z[24]);
endmodule

module CSA_23_5_26_0_25_000 (C, S, X, Y, Z);
  output [26:4] C;
  output [26:0] S;
  input [23:5] X;
  input [26:0] Y;
  input [25:3] Z;
  UBCON_2_0 U0 (S[2:0], Y[2:0]);
  PureCSHA_4_3 U1 (C[5:4], S[4:3], Z[4:3], Y[4:3]);
  PureCSA_23_5 U2 (C[24:6], S[23:5], X[23:5], Z[23:5], Y[23:5]);
  PureCSHA_25_24 U3 (C[26:25], S[25:24], Y[25:24], Z[25:24]);
  UB1DCON_26 U4 (S[26], Y[26]);
endmodule

module CSA_24_9_24_11_25000 (C, S, X, Y, Z);
  output [25:12] C;
  output [25:9] S;
  input [24:9] X;
  input [24:11] Y;
  input [25:12] Z;
  UBCON_10_9 U0 (S[10:9], X[10:9]);
  UBHA_11 U1 (C[12], S[11], Y[11], X[11]);
  PureCSA_24_12 U2 (C[25:13], S[24:12], Z[24:12], Y[24:12], X[24:12]);
  UB1DCON_25 U3 (S[25], Z[25]);
endmodule

module CSA_26_4_26_0_26_000 (C, S, X, Y, Z);
  output [27:5] C;
  output [26:0] S;
  input [26:4] X;
  input [26:0] Y;
  input [26:13] Z;
  UBCON_3_0 U0 (S[3:0], Y[3:0]);
  PureCSHA_12_4 U1 (C[13:5], S[12:4], X[12:4], Y[12:4]);
  PureCSA_26_13 U2 (C[27:14], S[26:13], Z[26:13], X[26:13], Y[26:13]);
endmodule

module MultUB_STD_OS_CSe000 (P, IN1, IN2);
  output [28:0] P;
  input [13:0] IN1;
  input [13:0] IN2;
  wire [13:0] PP0;
  wire [14:1] PP1;
  wire [23:10] PP10;
  wire [24:11] PP11;
  wire [25:12] PP12;
  wire [26:13] PP13;
  wire [15:2] PP2;
  wire [16:3] PP3;
  wire [17:4] PP4;
  wire [18:5] PP5;
  wire [19:6] PP6;
  wire [20:7] PP7;
  wire [21:8] PP8;
  wire [22:9] PP9;
  wire [27:5] S1;
  wire [26:0] S2;
  UBPPG_13_0_13_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, IN1, IN2);
  OSTR_13_0_14_1_15000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13);
  UBCSe_27_5_26_0 U2 (P, S1, S2);
endmodule

module OSBODY_13_0_14_1_000 (S0, S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13);
  output [26:4] S0;
  output [26:0] S1;
  output [26:13] S2;
  input [13:0] PP0;
  input [14:1] PP1;
  input [23:10] PP10;
  input [24:11] PP11;
  input [25:12] PP12;
  input [26:13] PP13;
  input [15:2] PP2;
  input [16:3] PP3;
  input [17:4] PP4;
  input [18:5] PP5;
  input [19:6] PP6;
  input [20:7] PP7;
  input [21:8] PP8;
  input [22:9] PP9;
  wire [23:5] W0;
  wire [26:0] W1;
  wire [25:3] W2;
  OSBODY_13_0_14_1_001 U0 (W0, W1, W2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12);
  OSCON_23_5_26_0_2000 U1 (S0, S1, S2, W0, W1, W2, PP13);
endmodule

module OSBODY_13_0_14_1_001 (S0, S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12);
  output [23:5] S0;
  output [26:0] S1;
  output [25:3] S2;
  input [13:0] PP0;
  input [14:1] PP1;
  input [23:10] PP10;
  input [24:11] PP11;
  input [25:12] PP12;
  input [15:2] PP2;
  input [16:3] PP3;
  input [17:4] PP4;
  input [18:5] PP5;
  input [19:6] PP6;
  input [20:7] PP7;
  input [21:8] PP8;
  input [22:9] PP9;
  wire [19:4] W0;
  wire [22:0] W1;
  wire [21:3] W2;
  wire [25:12] W3;
  wire [25:9] W4;
  OSBODY_13_0_14_1_002 U0 (W0, W1, W2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8);
  UBARYACC_22_9_23_000 U1 (W3, W4, PP9, PP10, PP11, PP12);
  OSCON_19_4_22_0_2000 U2 (S0, S1, S2, W0, W1, W2, W3, W4);
endmodule

module OSBODY_13_0_14_1_002 (S0, S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8);
  output [19:4] S0;
  output [22:0] S1;
  output [21:3] S2;
  input [13:0] PP0;
  input [14:1] PP1;
  input [15:2] PP2;
  input [16:3] PP3;
  input [17:4] PP4;
  input [18:5] PP5;
  input [19:6] PP6;
  input [20:7] PP7;
  input [21:8] PP8;
  wire [16:3] W0;
  wire [18:0] W1;
  wire [18:3] W2;
  wire [21:8] W3;
  wire [21:6] W4;
  OSBODY_13_0_14_1_003 U0 (W0, W1, W2, PP0, PP1, PP2, PP3, PP4, PP5);
  UBARYACC_19_6_20_000 U1 (W3, W4, PP6, PP7, PP8);
  OSCON_16_3_18_0_1000 U2 (S0, S1, S2, W0, W1, W2, W3, W4);
endmodule

module OSBODY_13_0_14_1_003 (S0, S1, S2, PP0, PP1, PP2, PP3, PP4, PP5);
  output [16:3] S0;
  output [18:0] S1;
  output [18:3] S2;
  input [13:0] PP0;
  input [14:1] PP1;
  input [15:2] PP2;
  input [16:3] PP3;
  input [17:4] PP4;
  input [18:5] PP5;
  wire [15:2] W0;
  wire [15:0] W1;
  wire [16:3] W2;
  wire [17:4] W3;
  wire [18:5] W4;
  OSBODY_13_0_14_1_004 U0 (W0, W1, W2, PP0, PP1, PP2, PP3);
  UBARYACC_17_4_18_000 U1 (W3, W4, PP4, PP5);
  OSCON_15_2_15_0_1000 U2 (S0, S1, S2, W0, W1, W2, W3, W4);
endmodule

module OSBODY_13_0_14_1_004 (S0, S1, S2, PP0, PP1, PP2, PP3);
  output [15:2] S0;
  output [15:0] S1;
  output [16:3] S2;
  input [13:0] PP0;
  input [14:1] PP1;
  input [15:2] PP2;
  input [16:3] PP3;
  CSA_13_0_14_1_15_000 U0 (S0, S1, PP0, PP1, PP2);
  UBCON_16_3 U1 (S2, PP3);
endmodule

module OSCON_15_2_15_0_1000 (S0, S1, S2, IN0, IN1, IN2, IN3, IN4);
  output [16:3] S0;
  output [18:0] S1;
  output [18:3] S2;
  input [15:2] IN0;
  input [15:0] IN1;
  input [16:3] IN2;
  input [17:4] IN3;
  input [18:5] IN4;
  wire [18:5] W;
  CSA_16_3_17_4_18_000 U0 (W, S2, IN2, IN3, IN4);
  CSA_15_2_15_0_18_000 U1 (S0, S1, IN0, IN1, W);
endmodule

module OSCON_16_3_18_0_1000 (S0, S1, S2, IN0, IN1, IN2, IN3, IN4);
  output [19:4] S0;
  output [22:0] S1;
  output [21:3] S2;
  input [16:3] IN0;
  input [18:0] IN1;
  input [18:3] IN2;
  input [21:8] IN3;
  input [21:6] IN4;
  wire [22:7] W;
  CSA_18_3_21_8_21_000 U0 (W, S2, IN2, IN3, IN4);
  CSA_16_3_18_0_22_000 U1 (S0, S1, IN0, IN1, W);
endmodule

module OSCON_19_4_22_0_2000 (S0, S1, S2, IN0, IN1, IN2, IN3, IN4);
  output [23:5] S0;
  output [26:0] S1;
  output [25:3] S2;
  input [19:4] IN0;
  input [22:0] IN1;
  input [21:3] IN2;
  input [25:12] IN3;
  input [25:9] IN4;
  wire [26:10] W;
  CSA_21_3_25_12_25000 U0 (W, S2, IN2, IN3, IN4);
  CSA_19_4_22_0_26_000 U1 (S0, S1, IN0, IN1, W);
endmodule

module OSCON_23_5_26_0_2000 (S0, S1, S2, IN0, IN1, IN2, IN3);
  output [26:4] S0;
  output [26:0] S1;
  output [26:13] S2;
  input [23:5] IN0;
  input [26:0] IN1;
  input [25:3] IN2;
  input [26:13] IN3;
  UBCON_26_13 U0 (S2, IN3);
  CSA_23_5_26_0_25_000 U1 (S0, S1, IN0, IN1, IN2);
endmodule

module OSTR_13_0_14_1_15000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13);
  output [27:5] S1;
  output [26:0] S2;
  input [13:0] PP0;
  input [14:1] PP1;
  input [23:10] PP10;
  input [24:11] PP11;
  input [25:12] PP12;
  input [26:13] PP13;
  input [15:2] PP2;
  input [16:3] PP3;
  input [17:4] PP4;
  input [18:5] PP5;
  input [19:6] PP6;
  input [20:7] PP7;
  input [21:8] PP8;
  input [22:9] PP9;
  wire [26:4] W0;
  wire [26:0] W1;
  wire [26:13] W2;
  OSBODY_13_0_14_1_000 U0 (W0, W1, W2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13);
  CSA_26_4_26_0_26_000 U1 (S1, S2, W0, W1, W2);
endmodule

module PureCSA_13_2 (C, S, X, Y, Z);
  output [14:3] C;
  output [13:2] S;
  input [13:2] X;
  input [13:2] Y;
  input [13:2] Z;
  UBFA_2 U0 (C[3], S[2], X[2], Y[2], Z[2]);
  UBFA_3 U1 (C[4], S[3], X[3], Y[3], Z[3]);
  UBFA_4 U2 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U3 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U4 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U5 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U6 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U7 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U8 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U9 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U10 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U11 (C[14], S[13], X[13], Y[13], Z[13]);
endmodule

module PureCSA_15_5 (C, S, X, Y, Z);
  output [16:6] C;
  output [15:5] S;
  input [15:5] X;
  input [15:5] Y;
  input [15:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U3 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U4 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U5 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U6 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U7 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U8 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U9 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U10 (C[16], S[15], X[15], Y[15], Z[15]);
endmodule

module PureCSA_16_5 (C, S, X, Y, Z);
  output [17:6] C;
  output [16:5] S;
  input [16:5] X;
  input [16:5] Y;
  input [16:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U3 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U4 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U5 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U6 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U7 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U8 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U9 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U10 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U11 (C[17], S[16], X[16], Y[16], Z[16]);
endmodule

module PureCSA_16_7 (C, S, X, Y, Z);
  output [17:8] C;
  output [16:7] S;
  input [16:7] X;
  input [16:7] Y;
  input [16:7] Z;
  UBFA_7 U0 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U1 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U2 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U3 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U4 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U5 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U6 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U7 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U8 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U9 (C[17], S[16], X[16], Y[16], Z[16]);
endmodule

module PureCSA_18_8 (C, S, X, Y, Z);
  output [19:9] C;
  output [18:8] S;
  input [18:8] X;
  input [18:8] Y;
  input [18:8] Z;
  UBFA_8 U0 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U1 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U2 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U3 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U4 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U5 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U6 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U7 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U8 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U9 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U10 (C[19], S[18], X[18], Y[18], Z[18]);
endmodule

module PureCSA_19_10 (C, S, X, Y, Z);
  output [20:11] C;
  output [19:10] S;
  input [19:10] X;
  input [19:10] Y;
  input [19:10] Z;
  UBFA_10 U0 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U1 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U2 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U3 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U4 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U5 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U6 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U7 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U8 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U9 (C[20], S[19], X[19], Y[19], Z[19]);
endmodule

module PureCSA_19_8 (C, S, X, Y, Z);
  output [20:9] C;
  output [19:8] S;
  input [19:8] X;
  input [19:8] Y;
  input [19:8] Z;
  UBFA_8 U0 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U1 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U2 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U3 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U4 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U5 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U6 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U7 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U8 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U9 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U10 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U11 (C[20], S[19], X[19], Y[19], Z[19]);
endmodule

module PureCSA_21_12 (C, S, X, Y, Z);
  output [22:13] C;
  output [21:12] S;
  input [21:12] X;
  input [21:12] Y;
  input [21:12] Z;
  UBFA_12 U0 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U1 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U2 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U3 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U4 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U5 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U6 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U7 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U8 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U9 (C[22], S[21], X[21], Y[21], Z[21]);
endmodule

module PureCSA_22_11 (C, S, X, Y, Z);
  output [23:12] C;
  output [22:11] S;
  input [22:11] X;
  input [22:11] Y;
  input [22:11] Z;
  UBFA_11 U0 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U1 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U2 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U3 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U4 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U5 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U6 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U7 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U8 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U9 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U10 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U11 (C[23], S[22], X[22], Y[22], Z[22]);
endmodule

module PureCSA_23_5 (C, S, X, Y, Z);
  output [24:6] C;
  output [23:5] S;
  input [23:5] X;
  input [23:5] Y;
  input [23:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U3 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U4 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U5 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U6 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U7 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U8 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U9 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U10 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U11 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U12 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U13 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U14 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U15 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U16 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U17 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U18 (C[24], S[23], X[23], Y[23], Z[23]);
endmodule

module PureCSA_24_12 (C, S, X, Y, Z);
  output [25:13] C;
  output [24:12] S;
  input [24:12] X;
  input [24:12] Y;
  input [24:12] Z;
  UBFA_12 U0 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U1 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U2 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U3 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U4 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U5 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U6 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U7 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U8 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U9 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U10 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U11 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U12 (C[25], S[24], X[24], Y[24], Z[24]);
endmodule

module PureCSA_26_13 (C, S, X, Y, Z);
  output [27:14] C;
  output [26:13] S;
  input [26:13] X;
  input [26:13] Y;
  input [26:13] Z;
  UBFA_13 U0 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U1 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U2 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U3 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U4 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U5 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U6 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U7 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U8 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U9 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U10 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U11 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U12 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U13 (C[27], S[26], X[26], Y[26], Z[26]);
endmodule

module PureCSHA_11_9 (C, S, X, Y);
  output [12:10] C;
  output [11:9] S;
  input [11:9] X;
  input [11:9] Y;
  UBHA_9 U0 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U1 (C[11], S[10], X[10], Y[10]);
  UBHA_11 U2 (C[12], S[11], X[11], Y[11]);
endmodule

module PureCSHA_12_4 (C, S, X, Y);
  output [13:5] C;
  output [12:4] S;
  input [12:4] X;
  input [12:4] Y;
  UBHA_4 U0 (C[5], S[4], X[4], Y[4]);
  UBHA_5 U1 (C[6], S[5], X[5], Y[5]);
  UBHA_6 U2 (C[7], S[6], X[6], Y[6]);
  UBHA_7 U3 (C[8], S[7], X[7], Y[7]);
  UBHA_8 U4 (C[9], S[8], X[8], Y[8]);
  UBHA_9 U5 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U6 (C[11], S[10], X[10], Y[10]);
  UBHA_11 U7 (C[12], S[11], X[11], Y[11]);
  UBHA_12 U8 (C[13], S[12], X[12], Y[12]);
endmodule

module PureCSHA_18_17 (C, S, X, Y);
  output [19:18] C;
  output [18:17] S;
  input [18:17] X;
  input [18:17] Y;
  UBHA_17 U0 (C[18], S[17], X[17], Y[17]);
  UBHA_18 U1 (C[19], S[18], X[18], Y[18]);
endmodule

module PureCSHA_21_19 (C, S, X, Y);
  output [22:20] C;
  output [21:19] S;
  input [21:19] X;
  input [21:19] Y;
  UBHA_19 U0 (C[20], S[19], X[19], Y[19]);
  UBHA_20 U1 (C[21], S[20], X[20], Y[20]);
  UBHA_21 U2 (C[22], S[21], X[21], Y[21]);
endmodule

module PureCSHA_22_20 (C, S, X, Y);
  output [23:21] C;
  output [22:20] S;
  input [22:20] X;
  input [22:20] Y;
  UBHA_20 U0 (C[21], S[20], X[20], Y[20]);
  UBHA_21 U1 (C[22], S[21], X[21], Y[21]);
  UBHA_22 U2 (C[23], S[22], X[22], Y[22]);
endmodule

module PureCSHA_25_22 (C, S, X, Y);
  output [26:23] C;
  output [25:22] S;
  input [25:22] X;
  input [25:22] Y;
  UBHA_22 U0 (C[23], S[22], X[22], Y[22]);
  UBHA_23 U1 (C[24], S[23], X[23], Y[23]);
  UBHA_24 U2 (C[25], S[24], X[24], Y[24]);
  UBHA_25 U3 (C[26], S[25], X[25], Y[25]);
endmodule

module PureCSHA_25_24 (C, S, X, Y);
  output [26:25] C;
  output [25:24] S;
  input [25:24] X;
  input [25:24] Y;
  UBHA_24 U0 (C[25], S[24], X[24], Y[24]);
  UBHA_25 U1 (C[26], S[25], X[25], Y[25]);
endmodule

module PureCSHA_4_2 (C, S, X, Y);
  output [5:3] C;
  output [4:2] S;
  input [4:2] X;
  input [4:2] Y;
  UBHA_2 U0 (C[3], S[2], X[2], Y[2]);
  UBHA_3 U1 (C[4], S[3], X[3], Y[3]);
  UBHA_4 U2 (C[5], S[4], X[4], Y[4]);
endmodule

module PureCSHA_4_3 (C, S, X, Y);
  output [5:4] C;
  output [4:3] S;
  input [4:3] X;
  input [4:3] Y;
  UBHA_3 U0 (C[4], S[3], X[3], Y[3]);
  UBHA_4 U1 (C[5], S[4], X[4], Y[4]);
endmodule

module PureCSHA_6_3 (C, S, X, Y);
  output [7:4] C;
  output [6:3] S;
  input [6:3] X;
  input [6:3] Y;
  UBHA_3 U0 (C[4], S[3], X[3], Y[3]);
  UBHA_4 U1 (C[5], S[4], X[4], Y[4]);
  UBHA_5 U2 (C[6], S[5], X[5], Y[5]);
  UBHA_6 U3 (C[7], S[6], X[6], Y[6]);
endmodule

module PureCSHA_7_6 (C, S, X, Y);
  output [8:7] C;
  output [7:6] S;
  input [7:6] X;
  input [7:6] Y;
  UBHA_6 U0 (C[7], S[6], X[6], Y[6]);
  UBHA_7 U1 (C[8], S[7], X[7], Y[7]);
endmodule

module PureCSHA_9_4 (C, S, X, Y);
  output [10:5] C;
  output [9:4] S;
  input [9:4] X;
  input [9:4] Y;
  UBHA_4 U0 (C[5], S[4], X[4], Y[4]);
  UBHA_5 U1 (C[6], S[5], X[5], Y[5]);
  UBHA_6 U2 (C[7], S[6], X[6], Y[6]);
  UBHA_7 U3 (C[8], S[7], X[7], Y[7]);
  UBHA_8 U4 (C[9], S[8], X[8], Y[8]);
  UBHA_9 U5 (C[10], S[9], X[9], Y[9]);
endmodule

module UBARYACC_17_4_18_000 (S1, S2, PP0, PP1);
  output [17:4] S1;
  output [18:5] S2;
  input [17:4] PP0;
  input [18:5] PP1;
  UBCON_17_4 U0 (S1, PP0);
  UBCON_18_5 U1 (S2, PP1);
endmodule

module UBARYACC_19_6_20_000 (S1, S2, PP0, PP1, PP2);
  output [21:8] S1;
  output [21:6] S2;
  input [19:6] PP0;
  input [20:7] PP1;
  input [21:8] PP2;
  CSA_19_6_20_7_21_000 U0 (S1, S2, PP0, PP1, PP2);
endmodule

module UBARYACC_22_9_23_000 (S1, S2, PP0, PP1, PP2, PP3);
  output [25:12] S1;
  output [25:9] S2;
  input [22:9] PP0;
  input [23:10] PP1;
  input [24:11] PP2;
  input [25:12] PP3;
  wire [24:11] IC0;
  wire [24:9] IS0;
  CSA_22_9_23_10_24000 U0 (IC0, IS0, PP0, PP1, PP2);
  CSA_24_9_24_11_25000 U1 (S1, S2, IS0, IC0, PP3);
endmodule

module UBCON_10_9 (O, I);
  output [10:9] O;
  input [10:9] I;
  UB1DCON_9 U0 (O[9], I[9]);
  UB1DCON_10 U1 (O[10], I[10]);
endmodule

module UBCON_16_3 (O, I);
  output [16:3] O;
  input [16:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
  UB1DCON_6 U3 (O[6], I[6]);
  UB1DCON_7 U4 (O[7], I[7]);
  UB1DCON_8 U5 (O[8], I[8]);
  UB1DCON_9 U6 (O[9], I[9]);
  UB1DCON_10 U7 (O[10], I[10]);
  UB1DCON_11 U8 (O[11], I[11]);
  UB1DCON_12 U9 (O[12], I[12]);
  UB1DCON_13 U10 (O[13], I[13]);
  UB1DCON_14 U11 (O[14], I[14]);
  UB1DCON_15 U12 (O[15], I[15]);
  UB1DCON_16 U13 (O[16], I[16]);
endmodule

module UBCON_17_4 (O, I);
  output [17:4] O;
  input [17:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
  UB1DCON_11 U7 (O[11], I[11]);
  UB1DCON_12 U8 (O[12], I[12]);
  UB1DCON_13 U9 (O[13], I[13]);
  UB1DCON_14 U10 (O[14], I[14]);
  UB1DCON_15 U11 (O[15], I[15]);
  UB1DCON_16 U12 (O[16], I[16]);
  UB1DCON_17 U13 (O[17], I[17]);
endmodule

module UBCON_18_16 (O, I);
  output [18:16] O;
  input [18:16] I;
  UB1DCON_16 U0 (O[16], I[16]);
  UB1DCON_17 U1 (O[17], I[17]);
  UB1DCON_18 U2 (O[18], I[18]);
endmodule

module UBCON_18_5 (O, I);
  output [18:5] O;
  input [18:5] I;
  UB1DCON_5 U0 (O[5], I[5]);
  UB1DCON_6 U1 (O[6], I[6]);
  UB1DCON_7 U2 (O[7], I[7]);
  UB1DCON_8 U3 (O[8], I[8]);
  UB1DCON_9 U4 (O[9], I[9]);
  UB1DCON_10 U5 (O[10], I[10]);
  UB1DCON_11 U6 (O[11], I[11]);
  UB1DCON_12 U7 (O[12], I[12]);
  UB1DCON_13 U8 (O[13], I[13]);
  UB1DCON_14 U9 (O[14], I[14]);
  UB1DCON_15 U10 (O[15], I[15]);
  UB1DCON_16 U11 (O[16], I[16]);
  UB1DCON_17 U12 (O[17], I[17]);
  UB1DCON_18 U13 (O[18], I[18]);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_22_19 (O, I);
  output [22:19] O;
  input [22:19] I;
  UB1DCON_19 U0 (O[19], I[19]);
  UB1DCON_20 U1 (O[20], I[20]);
  UB1DCON_21 U2 (O[21], I[21]);
  UB1DCON_22 U3 (O[22], I[22]);
endmodule

module UBCON_26_13 (O, I);
  output [26:13] O;
  input [26:13] I;
  UB1DCON_13 U0 (O[13], I[13]);
  UB1DCON_14 U1 (O[14], I[14]);
  UB1DCON_15 U2 (O[15], I[15]);
  UB1DCON_16 U3 (O[16], I[16]);
  UB1DCON_17 U4 (O[17], I[17]);
  UB1DCON_18 U5 (O[18], I[18]);
  UB1DCON_19 U6 (O[19], I[19]);
  UB1DCON_20 U7 (O[20], I[20]);
  UB1DCON_21 U8 (O[21], I[21]);
  UB1DCON_22 U9 (O[22], I[22]);
  UB1DCON_23 U10 (O[23], I[23]);
  UB1DCON_24 U11 (O[24], I[24]);
  UB1DCON_25 U12 (O[25], I[25]);
  UB1DCON_26 U13 (O[26], I[26]);
endmodule

module UBCON_26_23 (O, I);
  output [26:23] O;
  input [26:23] I;
  UB1DCON_23 U0 (O[23], I[23]);
  UB1DCON_24 U1 (O[24], I[24]);
  UB1DCON_25 U2 (O[25], I[25]);
  UB1DCON_26 U3 (O[26], I[26]);
endmodule

module UBCON_26_5 (O, I);
  output [26:5] O;
  input [26:5] I;
  UB1DCON_5 U0 (O[5], I[5]);
  UB1DCON_6 U1 (O[6], I[6]);
  UB1DCON_7 U2 (O[7], I[7]);
  UB1DCON_8 U3 (O[8], I[8]);
  UB1DCON_9 U4 (O[9], I[9]);
  UB1DCON_10 U5 (O[10], I[10]);
  UB1DCON_11 U6 (O[11], I[11]);
  UB1DCON_12 U7 (O[12], I[12]);
  UB1DCON_13 U8 (O[13], I[13]);
  UB1DCON_14 U9 (O[14], I[14]);
  UB1DCON_15 U10 (O[15], I[15]);
  UB1DCON_16 U11 (O[16], I[16]);
  UB1DCON_17 U12 (O[17], I[17]);
  UB1DCON_18 U13 (O[18], I[18]);
  UB1DCON_19 U14 (O[19], I[19]);
  UB1DCON_20 U15 (O[20], I[20]);
  UB1DCON_21 U16 (O[21], I[21]);
  UB1DCON_22 U17 (O[22], I[22]);
  UB1DCON_23 U18 (O[23], I[23]);
  UB1DCON_24 U19 (O[24], I[24]);
  UB1DCON_25 U20 (O[25], I[25]);
  UB1DCON_26 U21 (O[26], I[26]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBCON_3_0 (O, I);
  output [3:0] O;
  input [3:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
endmodule

module UBCON_4_0 (O, I);
  output [4:0] O;
  input [4:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
endmodule

module UBCON_5_3 (O, I);
  output [5:3] O;
  input [5:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
endmodule

module UBCON_8_3 (O, I);
  output [8:3] O;
  input [8:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
  UB1DCON_6 U3 (O[6], I[6]);
  UB1DCON_7 U4 (O[7], I[7]);
  UB1DCON_8 U5 (O[8], I[8]);
endmodule

module UBCSe_27_5_26_0 (S, X, Y);
  output [28:0] S;
  input [27:5] X;
  input [26:0] Y;
  wire [27:5] Z;
  UBExtender_26_5_2000 U0 (Z[27:5], Y[26:5]);
  UBPureCSe_27_5 U1 (S[28:5], X[27:5], Z[27:5]);
  UBCON_4_0 U2 (S[4:0], Y[4:0]);
endmodule

module UBExtender_26_5_2000 (O, I);
  output [27:5] O;
  input [26:5] I;
  UBCON_26_5 U0 (O[26:5], I[26:5]);
  UBZero_27_27 U1 (O[27]);
endmodule

module UBPPG_13_0_13_0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, IN1, IN2);
  output [13:0] PP0;
  output [14:1] PP1;
  output [23:10] PP10;
  output [24:11] PP11;
  output [25:12] PP12;
  output [26:13] PP13;
  output [15:2] PP2;
  output [16:3] PP3;
  output [17:4] PP4;
  output [18:5] PP5;
  output [19:6] PP6;
  output [20:7] PP7;
  output [21:8] PP8;
  output [22:9] PP9;
  input [13:0] IN1;
  input [13:0] IN2;
  UBVPPG_13_0_0 U0 (PP0, IN1, IN2[0]);
  UBVPPG_13_0_1 U1 (PP1, IN1, IN2[1]);
  UBVPPG_13_0_2 U2 (PP2, IN1, IN2[2]);
  UBVPPG_13_0_3 U3 (PP3, IN1, IN2[3]);
  UBVPPG_13_0_4 U4 (PP4, IN1, IN2[4]);
  UBVPPG_13_0_5 U5 (PP5, IN1, IN2[5]);
  UBVPPG_13_0_6 U6 (PP6, IN1, IN2[6]);
  UBVPPG_13_0_7 U7 (PP7, IN1, IN2[7]);
  UBVPPG_13_0_8 U8 (PP8, IN1, IN2[8]);
  UBVPPG_13_0_9 U9 (PP9, IN1, IN2[9]);
  UBVPPG_13_0_10 U10 (PP10, IN1, IN2[10]);
  UBVPPG_13_0_11 U11 (PP11, IN1, IN2[11]);
  UBVPPG_13_0_12 U12 (PP12, IN1, IN2[12]);
  UBVPPG_13_0_13 U13 (PP13, IN1, IN2[13]);
endmodule

module UBPureCSe_27_5 (S, X, Y);
  output [28:5] S;
  input [27:5] X;
  input [27:5] Y;
  wire C;
  UBPriCSlA_27_5 U0 (S, X, Y, C);
  UBZero_5_5 U1 (C);
endmodule

module UBRCB_11_9 (Co, S, X, Y, Ci);
  output Co;
  output [11:9] S;
  input Ci;
  input [11:9] X;
  input [11:9] Y;
  wire C10;
  wire C11;
  UBFA_9 U0 (C10, S[9], X[9], Y[9], Ci);
  UBFA_10 U1 (C11, S[10], X[10], Y[10], C10);
  UBFA_11 U2 (Co, S[11], X[11], Y[11], C11);
endmodule

module UBRCB_15_12 (Co, S, X, Y, Ci);
  output Co;
  output [15:12] S;
  input Ci;
  input [15:12] X;
  input [15:12] Y;
  wire C13;
  wire C14;
  wire C15;
  UBFA_12 U0 (C13, S[12], X[12], Y[12], Ci);
  UBFA_13 U1 (C14, S[13], X[13], Y[13], C13);
  UBFA_14 U2 (C15, S[14], X[14], Y[14], C14);
  UBFA_15 U3 (Co, S[15], X[15], Y[15], C15);
endmodule

module UBRCB_20_16 (Co, S, X, Y, Ci);
  output Co;
  output [20:16] S;
  input Ci;
  input [20:16] X;
  input [20:16] Y;
  wire C17;
  wire C18;
  wire C19;
  wire C20;
  UBFA_16 U0 (C17, S[16], X[16], Y[16], Ci);
  UBFA_17 U1 (C18, S[17], X[17], Y[17], C17);
  UBFA_18 U2 (C19, S[18], X[18], Y[18], C18);
  UBFA_19 U3 (C20, S[19], X[19], Y[19], C19);
  UBFA_20 U4 (Co, S[20], X[20], Y[20], C20);
endmodule

module UBRCB_26_21 (Co, S, X, Y, Ci);
  output Co;
  output [26:21] S;
  input Ci;
  input [26:21] X;
  input [26:21] Y;
  wire C22;
  wire C23;
  wire C24;
  wire C25;
  wire C26;
  UBFA_21 U0 (C22, S[21], X[21], Y[21], Ci);
  UBFA_22 U1 (C23, S[22], X[22], Y[22], C22);
  UBFA_23 U2 (C24, S[23], X[23], Y[23], C23);
  UBFA_24 U3 (C25, S[24], X[24], Y[24], C24);
  UBFA_25 U4 (C26, S[25], X[25], Y[25], C25);
  UBFA_26 U5 (Co, S[26], X[26], Y[26], C26);
endmodule

module UBRCB_27_27 (Co, S, X, Y, Ci);
  output Co;
  output S;
  input Ci;
  input X;
  input Y;
  UBFA_27 U0 (Co, S, X, Y, Ci);
endmodule

module UBRCB_5_5 (Co, S, X, Y, Ci);
  output Co;
  output S;
  input Ci;
  input X;
  input Y;
  UBFA_5 U0 (Co, S, X, Y, Ci);
endmodule

module UBRCB_6_6 (Co, S, X, Y, Ci);
  output Co;
  output S;
  input Ci;
  input X;
  input Y;
  UBFA_6 U0 (Co, S, X, Y, Ci);
endmodule

module UBRCB_8_7 (Co, S, X, Y, Ci);
  output Co;
  output [8:7] S;
  input Ci;
  input [8:7] X;
  input [8:7] Y;
  wire C8;
  UBFA_7 U0 (C8, S[7], X[7], Y[7], Ci);
  UBFA_8 U1 (Co, S[8], X[8], Y[8], C8);
endmodule

module UBVPPG_13_0_0 (O, IN1, IN2);
  output [13:0] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
  UB1BPPG_6_0 U6 (O[6], IN1[6], IN2);
  UB1BPPG_7_0 U7 (O[7], IN1[7], IN2);
  UB1BPPG_8_0 U8 (O[8], IN1[8], IN2);
  UB1BPPG_9_0 U9 (O[9], IN1[9], IN2);
  UB1BPPG_10_0 U10 (O[10], IN1[10], IN2);
  UB1BPPG_11_0 U11 (O[11], IN1[11], IN2);
  UB1BPPG_12_0 U12 (O[12], IN1[12], IN2);
  UB1BPPG_13_0 U13 (O[13], IN1[13], IN2);
endmodule

module UBVPPG_13_0_1 (O, IN1, IN2);
  output [14:1] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_1 U0 (O[1], IN1[0], IN2);
  UB1BPPG_1_1 U1 (O[2], IN1[1], IN2);
  UB1BPPG_2_1 U2 (O[3], IN1[2], IN2);
  UB1BPPG_3_1 U3 (O[4], IN1[3], IN2);
  UB1BPPG_4_1 U4 (O[5], IN1[4], IN2);
  UB1BPPG_5_1 U5 (O[6], IN1[5], IN2);
  UB1BPPG_6_1 U6 (O[7], IN1[6], IN2);
  UB1BPPG_7_1 U7 (O[8], IN1[7], IN2);
  UB1BPPG_8_1 U8 (O[9], IN1[8], IN2);
  UB1BPPG_9_1 U9 (O[10], IN1[9], IN2);
  UB1BPPG_10_1 U10 (O[11], IN1[10], IN2);
  UB1BPPG_11_1 U11 (O[12], IN1[11], IN2);
  UB1BPPG_12_1 U12 (O[13], IN1[12], IN2);
  UB1BPPG_13_1 U13 (O[14], IN1[13], IN2);
endmodule

module UBVPPG_13_0_10 (O, IN1, IN2);
  output [23:10] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_10 U0 (O[10], IN1[0], IN2);
  UB1BPPG_1_10 U1 (O[11], IN1[1], IN2);
  UB1BPPG_2_10 U2 (O[12], IN1[2], IN2);
  UB1BPPG_3_10 U3 (O[13], IN1[3], IN2);
  UB1BPPG_4_10 U4 (O[14], IN1[4], IN2);
  UB1BPPG_5_10 U5 (O[15], IN1[5], IN2);
  UB1BPPG_6_10 U6 (O[16], IN1[6], IN2);
  UB1BPPG_7_10 U7 (O[17], IN1[7], IN2);
  UB1BPPG_8_10 U8 (O[18], IN1[8], IN2);
  UB1BPPG_9_10 U9 (O[19], IN1[9], IN2);
  UB1BPPG_10_10 U10 (O[20], IN1[10], IN2);
  UB1BPPG_11_10 U11 (O[21], IN1[11], IN2);
  UB1BPPG_12_10 U12 (O[22], IN1[12], IN2);
  UB1BPPG_13_10 U13 (O[23], IN1[13], IN2);
endmodule

module UBVPPG_13_0_11 (O, IN1, IN2);
  output [24:11] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_11 U0 (O[11], IN1[0], IN2);
  UB1BPPG_1_11 U1 (O[12], IN1[1], IN2);
  UB1BPPG_2_11 U2 (O[13], IN1[2], IN2);
  UB1BPPG_3_11 U3 (O[14], IN1[3], IN2);
  UB1BPPG_4_11 U4 (O[15], IN1[4], IN2);
  UB1BPPG_5_11 U5 (O[16], IN1[5], IN2);
  UB1BPPG_6_11 U6 (O[17], IN1[6], IN2);
  UB1BPPG_7_11 U7 (O[18], IN1[7], IN2);
  UB1BPPG_8_11 U8 (O[19], IN1[8], IN2);
  UB1BPPG_9_11 U9 (O[20], IN1[9], IN2);
  UB1BPPG_10_11 U10 (O[21], IN1[10], IN2);
  UB1BPPG_11_11 U11 (O[22], IN1[11], IN2);
  UB1BPPG_12_11 U12 (O[23], IN1[12], IN2);
  UB1BPPG_13_11 U13 (O[24], IN1[13], IN2);
endmodule

module UBVPPG_13_0_12 (O, IN1, IN2);
  output [25:12] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_12 U0 (O[12], IN1[0], IN2);
  UB1BPPG_1_12 U1 (O[13], IN1[1], IN2);
  UB1BPPG_2_12 U2 (O[14], IN1[2], IN2);
  UB1BPPG_3_12 U3 (O[15], IN1[3], IN2);
  UB1BPPG_4_12 U4 (O[16], IN1[4], IN2);
  UB1BPPG_5_12 U5 (O[17], IN1[5], IN2);
  UB1BPPG_6_12 U6 (O[18], IN1[6], IN2);
  UB1BPPG_7_12 U7 (O[19], IN1[7], IN2);
  UB1BPPG_8_12 U8 (O[20], IN1[8], IN2);
  UB1BPPG_9_12 U9 (O[21], IN1[9], IN2);
  UB1BPPG_10_12 U10 (O[22], IN1[10], IN2);
  UB1BPPG_11_12 U11 (O[23], IN1[11], IN2);
  UB1BPPG_12_12 U12 (O[24], IN1[12], IN2);
  UB1BPPG_13_12 U13 (O[25], IN1[13], IN2);
endmodule

module UBVPPG_13_0_13 (O, IN1, IN2);
  output [26:13] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_13 U0 (O[13], IN1[0], IN2);
  UB1BPPG_1_13 U1 (O[14], IN1[1], IN2);
  UB1BPPG_2_13 U2 (O[15], IN1[2], IN2);
  UB1BPPG_3_13 U3 (O[16], IN1[3], IN2);
  UB1BPPG_4_13 U4 (O[17], IN1[4], IN2);
  UB1BPPG_5_13 U5 (O[18], IN1[5], IN2);
  UB1BPPG_6_13 U6 (O[19], IN1[6], IN2);
  UB1BPPG_7_13 U7 (O[20], IN1[7], IN2);
  UB1BPPG_8_13 U8 (O[21], IN1[8], IN2);
  UB1BPPG_9_13 U9 (O[22], IN1[9], IN2);
  UB1BPPG_10_13 U10 (O[23], IN1[10], IN2);
  UB1BPPG_11_13 U11 (O[24], IN1[11], IN2);
  UB1BPPG_12_13 U12 (O[25], IN1[12], IN2);
  UB1BPPG_13_13 U13 (O[26], IN1[13], IN2);
endmodule

module UBVPPG_13_0_2 (O, IN1, IN2);
  output [15:2] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
  UB1BPPG_6_2 U6 (O[8], IN1[6], IN2);
  UB1BPPG_7_2 U7 (O[9], IN1[7], IN2);
  UB1BPPG_8_2 U8 (O[10], IN1[8], IN2);
  UB1BPPG_9_2 U9 (O[11], IN1[9], IN2);
  UB1BPPG_10_2 U10 (O[12], IN1[10], IN2);
  UB1BPPG_11_2 U11 (O[13], IN1[11], IN2);
  UB1BPPG_12_2 U12 (O[14], IN1[12], IN2);
  UB1BPPG_13_2 U13 (O[15], IN1[13], IN2);
endmodule

module UBVPPG_13_0_3 (O, IN1, IN2);
  output [16:3] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_3 U0 (O[3], IN1[0], IN2);
  UB1BPPG_1_3 U1 (O[4], IN1[1], IN2);
  UB1BPPG_2_3 U2 (O[5], IN1[2], IN2);
  UB1BPPG_3_3 U3 (O[6], IN1[3], IN2);
  UB1BPPG_4_3 U4 (O[7], IN1[4], IN2);
  UB1BPPG_5_3 U5 (O[8], IN1[5], IN2);
  UB1BPPG_6_3 U6 (O[9], IN1[6], IN2);
  UB1BPPG_7_3 U7 (O[10], IN1[7], IN2);
  UB1BPPG_8_3 U8 (O[11], IN1[8], IN2);
  UB1BPPG_9_3 U9 (O[12], IN1[9], IN2);
  UB1BPPG_10_3 U10 (O[13], IN1[10], IN2);
  UB1BPPG_11_3 U11 (O[14], IN1[11], IN2);
  UB1BPPG_12_3 U12 (O[15], IN1[12], IN2);
  UB1BPPG_13_3 U13 (O[16], IN1[13], IN2);
endmodule

module UBVPPG_13_0_4 (O, IN1, IN2);
  output [17:4] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
  UB1BPPG_6_4 U6 (O[10], IN1[6], IN2);
  UB1BPPG_7_4 U7 (O[11], IN1[7], IN2);
  UB1BPPG_8_4 U8 (O[12], IN1[8], IN2);
  UB1BPPG_9_4 U9 (O[13], IN1[9], IN2);
  UB1BPPG_10_4 U10 (O[14], IN1[10], IN2);
  UB1BPPG_11_4 U11 (O[15], IN1[11], IN2);
  UB1BPPG_12_4 U12 (O[16], IN1[12], IN2);
  UB1BPPG_13_4 U13 (O[17], IN1[13], IN2);
endmodule

module UBVPPG_13_0_5 (O, IN1, IN2);
  output [18:5] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_5 U0 (O[5], IN1[0], IN2);
  UB1BPPG_1_5 U1 (O[6], IN1[1], IN2);
  UB1BPPG_2_5 U2 (O[7], IN1[2], IN2);
  UB1BPPG_3_5 U3 (O[8], IN1[3], IN2);
  UB1BPPG_4_5 U4 (O[9], IN1[4], IN2);
  UB1BPPG_5_5 U5 (O[10], IN1[5], IN2);
  UB1BPPG_6_5 U6 (O[11], IN1[6], IN2);
  UB1BPPG_7_5 U7 (O[12], IN1[7], IN2);
  UB1BPPG_8_5 U8 (O[13], IN1[8], IN2);
  UB1BPPG_9_5 U9 (O[14], IN1[9], IN2);
  UB1BPPG_10_5 U10 (O[15], IN1[10], IN2);
  UB1BPPG_11_5 U11 (O[16], IN1[11], IN2);
  UB1BPPG_12_5 U12 (O[17], IN1[12], IN2);
  UB1BPPG_13_5 U13 (O[18], IN1[13], IN2);
endmodule

module UBVPPG_13_0_6 (O, IN1, IN2);
  output [19:6] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_6 U0 (O[6], IN1[0], IN2);
  UB1BPPG_1_6 U1 (O[7], IN1[1], IN2);
  UB1BPPG_2_6 U2 (O[8], IN1[2], IN2);
  UB1BPPG_3_6 U3 (O[9], IN1[3], IN2);
  UB1BPPG_4_6 U4 (O[10], IN1[4], IN2);
  UB1BPPG_5_6 U5 (O[11], IN1[5], IN2);
  UB1BPPG_6_6 U6 (O[12], IN1[6], IN2);
  UB1BPPG_7_6 U7 (O[13], IN1[7], IN2);
  UB1BPPG_8_6 U8 (O[14], IN1[8], IN2);
  UB1BPPG_9_6 U9 (O[15], IN1[9], IN2);
  UB1BPPG_10_6 U10 (O[16], IN1[10], IN2);
  UB1BPPG_11_6 U11 (O[17], IN1[11], IN2);
  UB1BPPG_12_6 U12 (O[18], IN1[12], IN2);
  UB1BPPG_13_6 U13 (O[19], IN1[13], IN2);
endmodule

module UBVPPG_13_0_7 (O, IN1, IN2);
  output [20:7] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_7 U0 (O[7], IN1[0], IN2);
  UB1BPPG_1_7 U1 (O[8], IN1[1], IN2);
  UB1BPPG_2_7 U2 (O[9], IN1[2], IN2);
  UB1BPPG_3_7 U3 (O[10], IN1[3], IN2);
  UB1BPPG_4_7 U4 (O[11], IN1[4], IN2);
  UB1BPPG_5_7 U5 (O[12], IN1[5], IN2);
  UB1BPPG_6_7 U6 (O[13], IN1[6], IN2);
  UB1BPPG_7_7 U7 (O[14], IN1[7], IN2);
  UB1BPPG_8_7 U8 (O[15], IN1[8], IN2);
  UB1BPPG_9_7 U9 (O[16], IN1[9], IN2);
  UB1BPPG_10_7 U10 (O[17], IN1[10], IN2);
  UB1BPPG_11_7 U11 (O[18], IN1[11], IN2);
  UB1BPPG_12_7 U12 (O[19], IN1[12], IN2);
  UB1BPPG_13_7 U13 (O[20], IN1[13], IN2);
endmodule

module UBVPPG_13_0_8 (O, IN1, IN2);
  output [21:8] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_8 U0 (O[8], IN1[0], IN2);
  UB1BPPG_1_8 U1 (O[9], IN1[1], IN2);
  UB1BPPG_2_8 U2 (O[10], IN1[2], IN2);
  UB1BPPG_3_8 U3 (O[11], IN1[3], IN2);
  UB1BPPG_4_8 U4 (O[12], IN1[4], IN2);
  UB1BPPG_5_8 U5 (O[13], IN1[5], IN2);
  UB1BPPG_6_8 U6 (O[14], IN1[6], IN2);
  UB1BPPG_7_8 U7 (O[15], IN1[7], IN2);
  UB1BPPG_8_8 U8 (O[16], IN1[8], IN2);
  UB1BPPG_9_8 U9 (O[17], IN1[9], IN2);
  UB1BPPG_10_8 U10 (O[18], IN1[10], IN2);
  UB1BPPG_11_8 U11 (O[19], IN1[11], IN2);
  UB1BPPG_12_8 U12 (O[20], IN1[12], IN2);
  UB1BPPG_13_8 U13 (O[21], IN1[13], IN2);
endmodule

module UBVPPG_13_0_9 (O, IN1, IN2);
  output [22:9] O;
  input [13:0] IN1;
  input IN2;
  UB1BPPG_0_9 U0 (O[9], IN1[0], IN2);
  UB1BPPG_1_9 U1 (O[10], IN1[1], IN2);
  UB1BPPG_2_9 U2 (O[11], IN1[2], IN2);
  UB1BPPG_3_9 U3 (O[12], IN1[3], IN2);
  UB1BPPG_4_9 U4 (O[13], IN1[4], IN2);
  UB1BPPG_5_9 U5 (O[14], IN1[5], IN2);
  UB1BPPG_6_9 U6 (O[15], IN1[6], IN2);
  UB1BPPG_7_9 U7 (O[16], IN1[7], IN2);
  UB1BPPG_8_9 U8 (O[17], IN1[8], IN2);
  UB1BPPG_9_9 U9 (O[18], IN1[9], IN2);
  UB1BPPG_10_9 U10 (O[19], IN1[10], IN2);
  UB1BPPG_11_9 U11 (O[20], IN1[11], IN2);
  UB1BPPG_12_9 U12 (O[21], IN1[12], IN2);
  UB1BPPG_13_9 U13 (O[22], IN1[13], IN2);
endmodule

