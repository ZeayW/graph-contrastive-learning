/*----------------------------------------------------------------------------
  Copyright (c) 2019 Homma laboratory. All rights reserved.

  Top module: Multiplier_15_0_1000

  Number system: Unsigned binary
  Multiplicand length: 16
  Multiplier length: 16
  Partial product generation: Simple PPG
  Partial product accumulation: Dadda tree
  Final stage addition: Kogge-Stone adder
----------------------------------------------------------------------------*/

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_0_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UBHA_13(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_14(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBHA_14(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_15(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBHA_15(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_16(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBHA_16(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_17(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBFA_18(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_21(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_23(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_24(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_25(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_27(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_28(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_29(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_30(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_9(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBHA_10(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBHA_11(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_12(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBHA_12(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_13(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBFA_19(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBFA_20(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBFA_21(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBFA_22(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBHA_6(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBHA_7(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBHA_8(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBFA_23(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBFA_24(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBFA_25(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBHA_5(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBFA_26(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBFA_27(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBFA_28(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  GTECH_ADD_AB U0 (.A(X), .B(Y), .S(S), .COUT(C));
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module UBFA_29(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  GTECH_ADD_ABC U0 (.A(X), .B(Y), .C(Z), .S(S), .COUT(C));
endmodule

module GPGenerator(Go, Po, A, B);
  output Go;
  output Po;
  input A;
  input B;
  assign Go = A & B;
  assign Po = A ^ B;
endmodule

module CarryOperator(Go, Po, Gi1, Pi1, Gi2, Pi2);
  output Go;
  output Po;
  input Gi1;
  input Gi2;
  input Pi1;
  input Pi2;
  assign Go = Gi1 | ( Gi2 & Pi1 );
  assign Po = Pi1 & Pi2;
endmodule

module UBPriKSA_30_1(S, X, Y, Cin);
  output [31:1] S;
  input Cin;
  input [30:1] X;
  input [30:1] Y;
  wire [30:1] G0;
  wire [30:1] G1;
  wire [30:1] G2;
  wire [30:1] G3;
  wire [30:1] G4;
  wire [30:1] G5;
  wire [30:1] P0;
  wire [30:1] P1;
  wire [30:1] P2;
  wire [30:1] P3;
  wire [30:1] P4;
  wire [30:1] P5;
  assign P1[1] = P0[1];
  assign G1[1] = G0[1];
  assign P2[1] = P1[1];
  assign G2[1] = G1[1];
  assign P2[2] = P1[2];
  assign G2[2] = G1[2];
  assign P3[1] = P2[1];
  assign G3[1] = G2[1];
  assign P3[2] = P2[2];
  assign G3[2] = G2[2];
  assign P3[3] = P2[3];
  assign G3[3] = G2[3];
  assign P3[4] = P2[4];
  assign G3[4] = G2[4];
  assign P4[1] = P3[1];
  assign G4[1] = G3[1];
  assign P4[2] = P3[2];
  assign G4[2] = G3[2];
  assign P4[3] = P3[3];
  assign G4[3] = G3[3];
  assign P4[4] = P3[4];
  assign G4[4] = G3[4];
  assign P4[5] = P3[5];
  assign G4[5] = G3[5];
  assign P4[6] = P3[6];
  assign G4[6] = G3[6];
  assign P4[7] = P3[7];
  assign G4[7] = G3[7];
  assign P4[8] = P3[8];
  assign G4[8] = G3[8];
  assign P5[1] = P4[1];
  assign G5[1] = G4[1];
  assign P5[2] = P4[2];
  assign G5[2] = G4[2];
  assign P5[3] = P4[3];
  assign G5[3] = G4[3];
  assign P5[4] = P4[4];
  assign G5[4] = G4[4];
  assign P5[5] = P4[5];
  assign G5[5] = G4[5];
  assign P5[6] = P4[6];
  assign G5[6] = G4[6];
  assign P5[7] = P4[7];
  assign G5[7] = G4[7];
  assign P5[8] = P4[8];
  assign G5[8] = G4[8];
  assign P5[9] = P4[9];
  assign G5[9] = G4[9];
  assign P5[10] = P4[10];
  assign G5[10] = G4[10];
  assign P5[11] = P4[11];
  assign G5[11] = G4[11];
  assign P5[12] = P4[12];
  assign G5[12] = G4[12];
  assign P5[13] = P4[13];
  assign G5[13] = G4[13];
  assign P5[14] = P4[14];
  assign G5[14] = G4[14];
  assign P5[15] = P4[15];
  assign G5[15] = G4[15];
  assign P5[16] = P4[16];
  assign G5[16] = G4[16];
  assign S[1] = Cin ^ P0[1];
  assign S[2] = ( G5[1] | ( P5[1] & Cin ) ) ^ P0[2];
  assign S[3] = ( G5[2] | ( P5[2] & Cin ) ) ^ P0[3];
  assign S[4] = ( G5[3] | ( P5[3] & Cin ) ) ^ P0[4];
  assign S[5] = ( G5[4] | ( P5[4] & Cin ) ) ^ P0[5];
  assign S[6] = ( G5[5] | ( P5[5] & Cin ) ) ^ P0[6];
  assign S[7] = ( G5[6] | ( P5[6] & Cin ) ) ^ P0[7];
  assign S[8] = ( G5[7] | ( P5[7] & Cin ) ) ^ P0[8];
  assign S[9] = ( G5[8] | ( P5[8] & Cin ) ) ^ P0[9];
  assign S[10] = ( G5[9] | ( P5[9] & Cin ) ) ^ P0[10];
  assign S[11] = ( G5[10] | ( P5[10] & Cin ) ) ^ P0[11];
  assign S[12] = ( G5[11] | ( P5[11] & Cin ) ) ^ P0[12];
  assign S[13] = ( G5[12] | ( P5[12] & Cin ) ) ^ P0[13];
  assign S[14] = ( G5[13] | ( P5[13] & Cin ) ) ^ P0[14];
  assign S[15] = ( G5[14] | ( P5[14] & Cin ) ) ^ P0[15];
  assign S[16] = ( G5[15] | ( P5[15] & Cin ) ) ^ P0[16];
  assign S[17] = ( G5[16] | ( P5[16] & Cin ) ) ^ P0[17];
  assign S[18] = ( G5[17] | ( P5[17] & Cin ) ) ^ P0[18];
  assign S[19] = ( G5[18] | ( P5[18] & Cin ) ) ^ P0[19];
  assign S[20] = ( G5[19] | ( P5[19] & Cin ) ) ^ P0[20];
  assign S[21] = ( G5[20] | ( P5[20] & Cin ) ) ^ P0[21];
  assign S[22] = ( G5[21] | ( P5[21] & Cin ) ) ^ P0[22];
  assign S[23] = ( G5[22] | ( P5[22] & Cin ) ) ^ P0[23];
  assign S[24] = ( G5[23] | ( P5[23] & Cin ) ) ^ P0[24];
  assign S[25] = ( G5[24] | ( P5[24] & Cin ) ) ^ P0[25];
  assign S[26] = ( G5[25] | ( P5[25] & Cin ) ) ^ P0[26];
  assign S[27] = ( G5[26] | ( P5[26] & Cin ) ) ^ P0[27];
  assign S[28] = ( G5[27] | ( P5[27] & Cin ) ) ^ P0[28];
  assign S[29] = ( G5[28] | ( P5[28] & Cin ) ) ^ P0[29];
  assign S[30] = ( G5[29] | ( P5[29] & Cin ) ) ^ P0[30];
  assign S[31] = G5[30] | ( P5[30] & Cin );
  GPGenerator U0 (G0[1], P0[1], X[1], Y[1]);
  GPGenerator U1 (G0[2], P0[2], X[2], Y[2]);
  GPGenerator U2 (G0[3], P0[3], X[3], Y[3]);
  GPGenerator U3 (G0[4], P0[4], X[4], Y[4]);
  GPGenerator U4 (G0[5], P0[5], X[5], Y[5]);
  GPGenerator U5 (G0[6], P0[6], X[6], Y[6]);
  GPGenerator U6 (G0[7], P0[7], X[7], Y[7]);
  GPGenerator U7 (G0[8], P0[8], X[8], Y[8]);
  GPGenerator U8 (G0[9], P0[9], X[9], Y[9]);
  GPGenerator U9 (G0[10], P0[10], X[10], Y[10]);
  GPGenerator U10 (G0[11], P0[11], X[11], Y[11]);
  GPGenerator U11 (G0[12], P0[12], X[12], Y[12]);
  GPGenerator U12 (G0[13], P0[13], X[13], Y[13]);
  GPGenerator U13 (G0[14], P0[14], X[14], Y[14]);
  GPGenerator U14 (G0[15], P0[15], X[15], Y[15]);
  GPGenerator U15 (G0[16], P0[16], X[16], Y[16]);
  GPGenerator U16 (G0[17], P0[17], X[17], Y[17]);
  GPGenerator U17 (G0[18], P0[18], X[18], Y[18]);
  GPGenerator U18 (G0[19], P0[19], X[19], Y[19]);
  GPGenerator U19 (G0[20], P0[20], X[20], Y[20]);
  GPGenerator U20 (G0[21], P0[21], X[21], Y[21]);
  GPGenerator U21 (G0[22], P0[22], X[22], Y[22]);
  GPGenerator U22 (G0[23], P0[23], X[23], Y[23]);
  GPGenerator U23 (G0[24], P0[24], X[24], Y[24]);
  GPGenerator U24 (G0[25], P0[25], X[25], Y[25]);
  GPGenerator U25 (G0[26], P0[26], X[26], Y[26]);
  GPGenerator U26 (G0[27], P0[27], X[27], Y[27]);
  GPGenerator U27 (G0[28], P0[28], X[28], Y[28]);
  GPGenerator U28 (G0[29], P0[29], X[29], Y[29]);
  GPGenerator U29 (G0[30], P0[30], X[30], Y[30]);
  CarryOperator U30 (G1[2], P1[2], G0[2], P0[2], G0[1], P0[1]);
  CarryOperator U31 (G1[3], P1[3], G0[3], P0[3], G0[2], P0[2]);
  CarryOperator U32 (G1[4], P1[4], G0[4], P0[4], G0[3], P0[3]);
  CarryOperator U33 (G1[5], P1[5], G0[5], P0[5], G0[4], P0[4]);
  CarryOperator U34 (G1[6], P1[6], G0[6], P0[6], G0[5], P0[5]);
  CarryOperator U35 (G1[7], P1[7], G0[7], P0[7], G0[6], P0[6]);
  CarryOperator U36 (G1[8], P1[8], G0[8], P0[8], G0[7], P0[7]);
  CarryOperator U37 (G1[9], P1[9], G0[9], P0[9], G0[8], P0[8]);
  CarryOperator U38 (G1[10], P1[10], G0[10], P0[10], G0[9], P0[9]);
  CarryOperator U39 (G1[11], P1[11], G0[11], P0[11], G0[10], P0[10]);
  CarryOperator U40 (G1[12], P1[12], G0[12], P0[12], G0[11], P0[11]);
  CarryOperator U41 (G1[13], P1[13], G0[13], P0[13], G0[12], P0[12]);
  CarryOperator U42 (G1[14], P1[14], G0[14], P0[14], G0[13], P0[13]);
  CarryOperator U43 (G1[15], P1[15], G0[15], P0[15], G0[14], P0[14]);
  CarryOperator U44 (G1[16], P1[16], G0[16], P0[16], G0[15], P0[15]);
  CarryOperator U45 (G1[17], P1[17], G0[17], P0[17], G0[16], P0[16]);
  CarryOperator U46 (G1[18], P1[18], G0[18], P0[18], G0[17], P0[17]);
  CarryOperator U47 (G1[19], P1[19], G0[19], P0[19], G0[18], P0[18]);
  CarryOperator U48 (G1[20], P1[20], G0[20], P0[20], G0[19], P0[19]);
  CarryOperator U49 (G1[21], P1[21], G0[21], P0[21], G0[20], P0[20]);
  CarryOperator U50 (G1[22], P1[22], G0[22], P0[22], G0[21], P0[21]);
  CarryOperator U51 (G1[23], P1[23], G0[23], P0[23], G0[22], P0[22]);
  CarryOperator U52 (G1[24], P1[24], G0[24], P0[24], G0[23], P0[23]);
  CarryOperator U53 (G1[25], P1[25], G0[25], P0[25], G0[24], P0[24]);
  CarryOperator U54 (G1[26], P1[26], G0[26], P0[26], G0[25], P0[25]);
  CarryOperator U55 (G1[27], P1[27], G0[27], P0[27], G0[26], P0[26]);
  CarryOperator U56 (G1[28], P1[28], G0[28], P0[28], G0[27], P0[27]);
  CarryOperator U57 (G1[29], P1[29], G0[29], P0[29], G0[28], P0[28]);
  CarryOperator U58 (G1[30], P1[30], G0[30], P0[30], G0[29], P0[29]);
  CarryOperator U59 (G2[3], P2[3], G1[3], P1[3], G1[1], P1[1]);
  CarryOperator U60 (G2[4], P2[4], G1[4], P1[4], G1[2], P1[2]);
  CarryOperator U61 (G2[5], P2[5], G1[5], P1[5], G1[3], P1[3]);
  CarryOperator U62 (G2[6], P2[6], G1[6], P1[6], G1[4], P1[4]);
  CarryOperator U63 (G2[7], P2[7], G1[7], P1[7], G1[5], P1[5]);
  CarryOperator U64 (G2[8], P2[8], G1[8], P1[8], G1[6], P1[6]);
  CarryOperator U65 (G2[9], P2[9], G1[9], P1[9], G1[7], P1[7]);
  CarryOperator U66 (G2[10], P2[10], G1[10], P1[10], G1[8], P1[8]);
  CarryOperator U67 (G2[11], P2[11], G1[11], P1[11], G1[9], P1[9]);
  CarryOperator U68 (G2[12], P2[12], G1[12], P1[12], G1[10], P1[10]);
  CarryOperator U69 (G2[13], P2[13], G1[13], P1[13], G1[11], P1[11]);
  CarryOperator U70 (G2[14], P2[14], G1[14], P1[14], G1[12], P1[12]);
  CarryOperator U71 (G2[15], P2[15], G1[15], P1[15], G1[13], P1[13]);
  CarryOperator U72 (G2[16], P2[16], G1[16], P1[16], G1[14], P1[14]);
  CarryOperator U73 (G2[17], P2[17], G1[17], P1[17], G1[15], P1[15]);
  CarryOperator U74 (G2[18], P2[18], G1[18], P1[18], G1[16], P1[16]);
  CarryOperator U75 (G2[19], P2[19], G1[19], P1[19], G1[17], P1[17]);
  CarryOperator U76 (G2[20], P2[20], G1[20], P1[20], G1[18], P1[18]);
  CarryOperator U77 (G2[21], P2[21], G1[21], P1[21], G1[19], P1[19]);
  CarryOperator U78 (G2[22], P2[22], G1[22], P1[22], G1[20], P1[20]);
  CarryOperator U79 (G2[23], P2[23], G1[23], P1[23], G1[21], P1[21]);
  CarryOperator U80 (G2[24], P2[24], G1[24], P1[24], G1[22], P1[22]);
  CarryOperator U81 (G2[25], P2[25], G1[25], P1[25], G1[23], P1[23]);
  CarryOperator U82 (G2[26], P2[26], G1[26], P1[26], G1[24], P1[24]);
  CarryOperator U83 (G2[27], P2[27], G1[27], P1[27], G1[25], P1[25]);
  CarryOperator U84 (G2[28], P2[28], G1[28], P1[28], G1[26], P1[26]);
  CarryOperator U85 (G2[29], P2[29], G1[29], P1[29], G1[27], P1[27]);
  CarryOperator U86 (G2[30], P2[30], G1[30], P1[30], G1[28], P1[28]);
  CarryOperator U87 (G3[5], P3[5], G2[5], P2[5], G2[1], P2[1]);
  CarryOperator U88 (G3[6], P3[6], G2[6], P2[6], G2[2], P2[2]);
  CarryOperator U89 (G3[7], P3[7], G2[7], P2[7], G2[3], P2[3]);
  CarryOperator U90 (G3[8], P3[8], G2[8], P2[8], G2[4], P2[4]);
  CarryOperator U91 (G3[9], P3[9], G2[9], P2[9], G2[5], P2[5]);
  CarryOperator U92 (G3[10], P3[10], G2[10], P2[10], G2[6], P2[6]);
  CarryOperator U93 (G3[11], P3[11], G2[11], P2[11], G2[7], P2[7]);
  CarryOperator U94 (G3[12], P3[12], G2[12], P2[12], G2[8], P2[8]);
  CarryOperator U95 (G3[13], P3[13], G2[13], P2[13], G2[9], P2[9]);
  CarryOperator U96 (G3[14], P3[14], G2[14], P2[14], G2[10], P2[10]);
  CarryOperator U97 (G3[15], P3[15], G2[15], P2[15], G2[11], P2[11]);
  CarryOperator U98 (G3[16], P3[16], G2[16], P2[16], G2[12], P2[12]);
  CarryOperator U99 (G3[17], P3[17], G2[17], P2[17], G2[13], P2[13]);
  CarryOperator U100 (G3[18], P3[18], G2[18], P2[18], G2[14], P2[14]);
  CarryOperator U101 (G3[19], P3[19], G2[19], P2[19], G2[15], P2[15]);
  CarryOperator U102 (G3[20], P3[20], G2[20], P2[20], G2[16], P2[16]);
  CarryOperator U103 (G3[21], P3[21], G2[21], P2[21], G2[17], P2[17]);
  CarryOperator U104 (G3[22], P3[22], G2[22], P2[22], G2[18], P2[18]);
  CarryOperator U105 (G3[23], P3[23], G2[23], P2[23], G2[19], P2[19]);
  CarryOperator U106 (G3[24], P3[24], G2[24], P2[24], G2[20], P2[20]);
  CarryOperator U107 (G3[25], P3[25], G2[25], P2[25], G2[21], P2[21]);
  CarryOperator U108 (G3[26], P3[26], G2[26], P2[26], G2[22], P2[22]);
  CarryOperator U109 (G3[27], P3[27], G2[27], P2[27], G2[23], P2[23]);
  CarryOperator U110 (G3[28], P3[28], G2[28], P2[28], G2[24], P2[24]);
  CarryOperator U111 (G3[29], P3[29], G2[29], P2[29], G2[25], P2[25]);
  CarryOperator U112 (G3[30], P3[30], G2[30], P2[30], G2[26], P2[26]);
  CarryOperator U113 (G4[9], P4[9], G3[9], P3[9], G3[1], P3[1]);
  CarryOperator U114 (G4[10], P4[10], G3[10], P3[10], G3[2], P3[2]);
  CarryOperator U115 (G4[11], P4[11], G3[11], P3[11], G3[3], P3[3]);
  CarryOperator U116 (G4[12], P4[12], G3[12], P3[12], G3[4], P3[4]);
  CarryOperator U117 (G4[13], P4[13], G3[13], P3[13], G3[5], P3[5]);
  CarryOperator U118 (G4[14], P4[14], G3[14], P3[14], G3[6], P3[6]);
  CarryOperator U119 (G4[15], P4[15], G3[15], P3[15], G3[7], P3[7]);
  CarryOperator U120 (G4[16], P4[16], G3[16], P3[16], G3[8], P3[8]);
  CarryOperator U121 (G4[17], P4[17], G3[17], P3[17], G3[9], P3[9]);
  CarryOperator U122 (G4[18], P4[18], G3[18], P3[18], G3[10], P3[10]);
  CarryOperator U123 (G4[19], P4[19], G3[19], P3[19], G3[11], P3[11]);
  CarryOperator U124 (G4[20], P4[20], G3[20], P3[20], G3[12], P3[12]);
  CarryOperator U125 (G4[21], P4[21], G3[21], P3[21], G3[13], P3[13]);
  CarryOperator U126 (G4[22], P4[22], G3[22], P3[22], G3[14], P3[14]);
  CarryOperator U127 (G4[23], P4[23], G3[23], P3[23], G3[15], P3[15]);
  CarryOperator U128 (G4[24], P4[24], G3[24], P3[24], G3[16], P3[16]);
  CarryOperator U129 (G4[25], P4[25], G3[25], P3[25], G3[17], P3[17]);
  CarryOperator U130 (G4[26], P4[26], G3[26], P3[26], G3[18], P3[18]);
  CarryOperator U131 (G4[27], P4[27], G3[27], P3[27], G3[19], P3[19]);
  CarryOperator U132 (G4[28], P4[28], G3[28], P3[28], G3[20], P3[20]);
  CarryOperator U133 (G4[29], P4[29], G3[29], P3[29], G3[21], P3[21]);
  CarryOperator U134 (G4[30], P4[30], G3[30], P3[30], G3[22], P3[22]);
  CarryOperator U135 (G5[17], P5[17], G4[17], P4[17], G4[1], P4[1]);
  CarryOperator U136 (G5[18], P5[18], G4[18], P4[18], G4[2], P4[2]);
  CarryOperator U137 (G5[19], P5[19], G4[19], P4[19], G4[3], P4[3]);
  CarryOperator U138 (G5[20], P5[20], G4[20], P4[20], G4[4], P4[4]);
  CarryOperator U139 (G5[21], P5[21], G4[21], P4[21], G4[5], P4[5]);
  CarryOperator U140 (G5[22], P5[22], G4[22], P4[22], G4[6], P4[6]);
  CarryOperator U141 (G5[23], P5[23], G4[23], P4[23], G4[7], P4[7]);
  CarryOperator U142 (G5[24], P5[24], G4[24], P4[24], G4[8], P4[8]);
  CarryOperator U143 (G5[25], P5[25], G4[25], P4[25], G4[9], P4[9]);
  CarryOperator U144 (G5[26], P5[26], G4[26], P4[26], G4[10], P4[10]);
  CarryOperator U145 (G5[27], P5[27], G4[27], P4[27], G4[11], P4[11]);
  CarryOperator U146 (G5[28], P5[28], G4[28], P4[28], G4[12], P4[12]);
  CarryOperator U147 (G5[29], P5[29], G4[29], P4[29], G4[13], P4[13]);
  CarryOperator U148 (G5[30], P5[30], G4[30], P4[30], G4[14], P4[14]);
endmodule

module UBZero_1_1(O);
  output [1:1] O;
  assign O[1] = 0;
endmodule

module Multiplier_15_0_1000(P, IN1, IN2);
  output [31:0] P;
  input [15:0] IN1;
  input [15:0] IN2;
  wire [31:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  assign P[12] = W[12];
  assign P[13] = W[13];
  assign P[14] = W[14];
  assign P[15] = W[15];
  assign P[16] = W[16];
  assign P[17] = W[17];
  assign P[18] = W[18];
  assign P[19] = W[19];
  assign P[20] = W[20];
  assign P[21] = W[21];
  assign P[22] = W[22];
  assign P[23] = W[23];
  assign P[24] = W[24];
  assign P[25] = W[25];
  assign P[26] = W[26];
  assign P[27] = W[27];
  assign P[28] = W[28];
  assign P[29] = W[29];
  assign P[30] = W[30];
  assign P[31] = W[31];
  MultUB_STD_DAD_KS000 U0 (W, IN1, IN2);
endmodule

module DADTR_15_0_16_1_1000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15);
  output [30:0] S1;
  output [30:1] S2;
  input [15:0] PP0;
  input [16:1] PP1;
  input [25:10] PP10;
  input [26:11] PP11;
  input [27:12] PP12;
  input [28:13] PP13;
  input [29:14] PP14;
  input [30:15] PP15;
  input [17:2] PP2;
  input [18:3] PP3;
  input [19:4] PP4;
  input [20:5] PP5;
  input [21:6] PP6;
  input [22:7] PP7;
  input [23:8] PP8;
  input [24:9] PP9;
  wire [30:0] W0;
  wire [29:1] W1;
  wire [20:10] W10;
  wire [19:11] W11;
  wire [19:12] W12;
  wire [28:2] W2;
  wire [27:3] W3;
  wire [26:4] W4;
  wire [25:5] W5;
  wire [24:6] W6;
  wire [23:7] W7;
  wire [22:8] W8;
  wire [21:9] W9;
  UBHA_13 U0 (W10[14], W12[13], PP0[13], PP1[13]);
  UBFA_14 U1 (W8[15], W11[14], PP0[14], PP1[14], PP2[14]);
  UBHA_14 U2 (W9[15], W12[14], PP3[14], PP4[14]);
  UBFA_15 U3 (W7[16], W10[15], PP0[15], PP1[15], PP2[15]);
  UBFA_15 U4 (W8[16], W11[15], PP3[15], PP4[15], PP5[15]);
  UBHA_15 U5 (W9[16], W12[15], PP6[15], PP7[15]);
  UBFA_16 U6 (W8[17], W10[16], PP1[16], PP2[16], PP3[16]);
  UBFA_16 U7 (W9[17], W11[16], PP4[16], PP5[16], PP6[16]);
  UBHA_16 U8 (W10[17], W12[16], PP7[16], PP8[16]);
  UBFA_17 U9 (W10[18], W11[17], PP2[17], PP3[17], PP4[17]);
  UBFA_17 U10 (W11[18], W12[17], PP5[17], PP6[17], PP7[17]);
  UBFA_18 U11 (W12[19], W12[18], PP3[18], PP4[18], PP5[18]);
  UBCON_12_0 U12 (W0[12:0], PP0[12:0]);
  UB1DCON_13 U13 (W0[13], PP2[13]);
  UB1DCON_14 U14 (W0[14], PP5[14]);
  UB1DCON_15 U15 (W0[15], PP8[15]);
  UB1DCON_16 U16 (W0[16], PP9[16]);
  UB1DCON_17 U17 (W0[17], PP8[17]);
  UB1DCON_18 U18 (W0[18], PP6[18]);
  UB1DCON_19 U19 (W0[19], PP4[19]);
  UB1DCON_20 U20 (W0[20], PP5[20]);
  UB1DCON_21 U21 (W0[21], PP6[21]);
  UB1DCON_22 U22 (W0[22], PP7[22]);
  UB1DCON_23 U23 (W0[23], PP8[23]);
  UB1DCON_24 U24 (W0[24], PP9[24]);
  UB1DCON_25 U25 (W0[25], PP10[25]);
  UB1DCON_26 U26 (W0[26], PP11[26]);
  UB1DCON_27 U27 (W0[27], PP12[27]);
  UB1DCON_28 U28 (W0[28], PP13[28]);
  UB1DCON_29 U29 (W0[29], PP14[29]);
  UB1DCON_30 U30 (W0[30], PP15[30]);
  UBCON_12_1 U31 (W1[12:1], PP1[12:1]);
  UB1DCON_13 U32 (W1[13], PP3[13]);
  UB1DCON_14 U33 (W1[14], PP6[14]);
  UB1DCON_15 U34 (W1[15], PP9[15]);
  UB1DCON_16 U35 (W1[16], PP10[16]);
  UB1DCON_17 U36 (W1[17], PP9[17]);
  UB1DCON_18 U37 (W1[18], PP7[18]);
  UB1DCON_19 U38 (W1[19], PP5[19]);
  UB1DCON_20 U39 (W1[20], PP6[20]);
  UB1DCON_21 U40 (W1[21], PP7[21]);
  UB1DCON_22 U41 (W1[22], PP8[22]);
  UB1DCON_23 U42 (W1[23], PP9[23]);
  UB1DCON_24 U43 (W1[24], PP10[24]);
  UB1DCON_25 U44 (W1[25], PP11[25]);
  UB1DCON_26 U45 (W1[26], PP12[26]);
  UB1DCON_27 U46 (W1[27], PP13[27]);
  UB1DCON_28 U47 (W1[28], PP14[28]);
  UB1DCON_29 U48 (W1[29], PP15[29]);
  UBCON_12_2 U49 (W2[12:2], PP2[12:2]);
  UB1DCON_13 U50 (W2[13], PP4[13]);
  UB1DCON_14 U51 (W2[14], PP7[14]);
  UB1DCON_15 U52 (W2[15], PP10[15]);
  UB1DCON_16 U53 (W2[16], PP11[16]);
  UB1DCON_17 U54 (W2[17], PP10[17]);
  UB1DCON_18 U55 (W2[18], PP8[18]);
  UB1DCON_19 U56 (W2[19], PP6[19]);
  UB1DCON_20 U57 (W2[20], PP7[20]);
  UB1DCON_21 U58 (W2[21], PP8[21]);
  UB1DCON_22 U59 (W2[22], PP9[22]);
  UB1DCON_23 U60 (W2[23], PP10[23]);
  UB1DCON_24 U61 (W2[24], PP11[24]);
  UB1DCON_25 U62 (W2[25], PP12[25]);
  UB1DCON_26 U63 (W2[26], PP13[26]);
  UB1DCON_27 U64 (W2[27], PP14[27]);
  UB1DCON_28 U65 (W2[28], PP15[28]);
  UBCON_12_3 U66 (W3[12:3], PP3[12:3]);
  UB1DCON_13 U67 (W3[13], PP5[13]);
  UB1DCON_14 U68 (W3[14], PP8[14]);
  UB1DCON_15 U69 (W3[15], PP11[15]);
  UB1DCON_16 U70 (W3[16], PP12[16]);
  UB1DCON_17 U71 (W3[17], PP11[17]);
  UB1DCON_18 U72 (W3[18], PP9[18]);
  UB1DCON_19 U73 (W3[19], PP7[19]);
  UB1DCON_20 U74 (W3[20], PP8[20]);
  UB1DCON_21 U75 (W3[21], PP9[21]);
  UB1DCON_22 U76 (W3[22], PP10[22]);
  UB1DCON_23 U77 (W3[23], PP11[23]);
  UB1DCON_24 U78 (W3[24], PP12[24]);
  UB1DCON_25 U79 (W3[25], PP13[25]);
  UB1DCON_26 U80 (W3[26], PP14[26]);
  UB1DCON_27 U81 (W3[27], PP15[27]);
  UBCON_12_4 U82 (W4[12:4], PP4[12:4]);
  UB1DCON_13 U83 (W4[13], PP6[13]);
  UB1DCON_14 U84 (W4[14], PP9[14]);
  UB1DCON_15 U85 (W4[15], PP12[15]);
  UB1DCON_16 U86 (W4[16], PP13[16]);
  UB1DCON_17 U87 (W4[17], PP12[17]);
  UB1DCON_18 U88 (W4[18], PP10[18]);
  UB1DCON_19 U89 (W4[19], PP8[19]);
  UB1DCON_20 U90 (W4[20], PP9[20]);
  UB1DCON_21 U91 (W4[21], PP10[21]);
  UB1DCON_22 U92 (W4[22], PP11[22]);
  UB1DCON_23 U93 (W4[23], PP12[23]);
  UB1DCON_24 U94 (W4[24], PP13[24]);
  UB1DCON_25 U95 (W4[25], PP14[25]);
  UB1DCON_26 U96 (W4[26], PP15[26]);
  UBCON_12_5 U97 (W5[12:5], PP5[12:5]);
  UB1DCON_13 U98 (W5[13], PP7[13]);
  UB1DCON_14 U99 (W5[14], PP10[14]);
  UB1DCON_15 U100 (W5[15], PP13[15]);
  UB1DCON_16 U101 (W5[16], PP14[16]);
  UB1DCON_17 U102 (W5[17], PP13[17]);
  UB1DCON_18 U103 (W5[18], PP11[18]);
  UB1DCON_19 U104 (W5[19], PP9[19]);
  UB1DCON_20 U105 (W5[20], PP10[20]);
  UB1DCON_21 U106 (W5[21], PP11[21]);
  UB1DCON_22 U107 (W5[22], PP12[22]);
  UB1DCON_23 U108 (W5[23], PP13[23]);
  UB1DCON_24 U109 (W5[24], PP14[24]);
  UB1DCON_25 U110 (W5[25], PP15[25]);
  UBCON_12_6 U111 (W6[12:6], PP6[12:6]);
  UB1DCON_13 U112 (W6[13], PP8[13]);
  UB1DCON_14 U113 (W6[14], PP11[14]);
  UB1DCON_15 U114 (W6[15], PP14[15]);
  UB1DCON_16 U115 (W6[16], PP15[16]);
  UB1DCON_17 U116 (W6[17], PP14[17]);
  UB1DCON_18 U117 (W6[18], PP12[18]);
  UB1DCON_19 U118 (W6[19], PP10[19]);
  UB1DCON_20 U119 (W6[20], PP11[20]);
  UB1DCON_21 U120 (W6[21], PP12[21]);
  UB1DCON_22 U121 (W6[22], PP13[22]);
  UB1DCON_23 U122 (W6[23], PP14[23]);
  UB1DCON_24 U123 (W6[24], PP15[24]);
  UBCON_12_7 U124 (W7[12:7], PP7[12:7]);
  UB1DCON_13 U125 (W7[13], PP9[13]);
  UB1DCON_14 U126 (W7[14], PP12[14]);
  UB1DCON_15 U127 (W7[15], PP15[15]);
  UB1DCON_17 U128 (W7[17], PP15[17]);
  UB1DCON_18 U129 (W7[18], PP13[18]);
  UB1DCON_19 U130 (W7[19], PP11[19]);
  UB1DCON_20 U131 (W7[20], PP12[20]);
  UB1DCON_21 U132 (W7[21], PP13[21]);
  UB1DCON_22 U133 (W7[22], PP14[22]);
  UB1DCON_23 U134 (W7[23], PP15[23]);
  UBCON_12_8 U135 (W8[12:8], PP8[12:8]);
  UB1DCON_13 U136 (W8[13], PP10[13]);
  UB1DCON_14 U137 (W8[14], PP13[14]);
  UB1DCON_18 U138 (W8[18], PP14[18]);
  UB1DCON_19 U139 (W8[19], PP12[19]);
  UB1DCON_20 U140 (W8[20], PP13[20]);
  UB1DCON_21 U141 (W8[21], PP14[21]);
  UB1DCON_22 U142 (W8[22], PP15[22]);
  UBCON_12_9 U143 (W9[12:9], PP9[12:9]);
  UB1DCON_13 U144 (W9[13], PP11[13]);
  UB1DCON_14 U145 (W9[14], PP14[14]);
  UB1DCON_18 U146 (W9[18], PP15[18]);
  UB1DCON_19 U147 (W9[19], PP13[19]);
  UB1DCON_20 U148 (W9[20], PP14[20]);
  UB1DCON_21 U149 (W9[21], PP15[21]);
  UBCON_12_10 U150 (W10[12:10], PP10[12:10]);
  UB1DCON_13 U151 (W10[13], PP12[13]);
  UB1DCON_19 U152 (W10[19], PP14[19]);
  UB1DCON_20 U153 (W10[20], PP15[20]);
  UBCON_12_11 U154 (W11[12:11], PP11[12:11]);
  UB1DCON_13 U155 (W11[13], PP13[13]);
  UB1DCON_19 U156 (W11[19], PP15[19]);
  UB1DCON_12 U157 (W12[12], PP12[12]);
  DADTR_30_0_29_1_2000 U158 (S1, S2, W0, W1, W2, W3, W4, W5, W6, W7, W8, W9, W10, W11, W12);
endmodule

module DADTR_30_0_29_1_2000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12);
  output [30:0] S1;
  output [30:1] S2;
  input [30:0] PP0;
  input [29:1] PP1;
  input [20:10] PP10;
  input [19:11] PP11;
  input [19:12] PP12;
  input [28:2] PP2;
  input [27:3] PP3;
  input [26:4] PP4;
  input [25:5] PP5;
  input [24:6] PP6;
  input [23:7] PP7;
  input [22:8] PP8;
  input [21:9] PP9;
  wire [30:0] W0;
  wire [29:1] W1;
  wire [28:2] W2;
  wire [27:3] W3;
  wire [26:4] W4;
  wire [25:5] W5;
  wire [24:6] W6;
  wire [23:7] W7;
  wire [23:8] W8;
  UBHA_9 U0 (W6[10], W8[9], PP0[9], PP1[9]);
  UBFA_10 U1 (W4[11], W7[10], PP0[10], PP1[10], PP2[10]);
  UBHA_10 U2 (W5[11], W8[10], PP3[10], PP4[10]);
  UBFA_11 U3 (W2[12], W6[11], PP0[11], PP1[11], PP2[11]);
  UBFA_11 U4 (W3[12], W7[11], PP3[11], PP4[11], PP5[11]);
  UBHA_11 U5 (W4[12], W8[11], PP6[11], PP7[11]);
  UBFA_12 U6 (W1[13], W5[12], PP0[12], PP1[12], PP2[12]);
  UBFA_12 U7 (W2[13], W6[12], PP3[12], PP4[12], PP5[12]);
  UBFA_12 U8 (W3[13], W7[12], PP6[12], PP7[12], PP8[12]);
  UBHA_12 U9 (W4[13], W8[12], PP9[12], PP10[12]);
  UBFA_13 U10 (W1[14], W5[13], PP0[13], PP1[13], PP2[13]);
  UBFA_13 U11 (W2[14], W6[13], PP3[13], PP4[13], PP5[13]);
  UBFA_13 U12 (W3[14], W7[13], PP6[13], PP7[13], PP8[13]);
  UBFA_13 U13 (W4[14], W8[13], PP9[13], PP10[13], PP11[13]);
  UBFA_14 U14 (W1[15], W5[14], PP0[14], PP1[14], PP2[14]);
  UBFA_14 U15 (W2[15], W6[14], PP3[14], PP4[14], PP5[14]);
  UBFA_14 U16 (W3[15], W7[14], PP6[14], PP7[14], PP8[14]);
  UBFA_14 U17 (W4[15], W8[14], PP9[14], PP10[14], PP11[14]);
  UBFA_15 U18 (W1[16], W5[15], PP0[15], PP1[15], PP2[15]);
  UBFA_15 U19 (W2[16], W6[15], PP3[15], PP4[15], PP5[15]);
  UBFA_15 U20 (W3[16], W7[15], PP6[15], PP7[15], PP8[15]);
  UBFA_15 U21 (W4[16], W8[15], PP9[15], PP10[15], PP11[15]);
  UBFA_16 U22 (W1[17], W5[16], PP0[16], PP1[16], PP2[16]);
  UBFA_16 U23 (W2[17], W6[16], PP3[16], PP4[16], PP5[16]);
  UBFA_16 U24 (W3[17], W7[16], PP6[16], PP7[16], PP8[16]);
  UBFA_16 U25 (W4[17], W8[16], PP9[16], PP10[16], PP11[16]);
  UBFA_17 U26 (W1[18], W5[17], PP0[17], PP1[17], PP2[17]);
  UBFA_17 U27 (W2[18], W6[17], PP3[17], PP4[17], PP5[17]);
  UBFA_17 U28 (W3[18], W7[17], PP6[17], PP7[17], PP8[17]);
  UBFA_17 U29 (W4[18], W8[17], PP9[17], PP10[17], PP11[17]);
  UBFA_18 U30 (W1[19], W5[18], PP0[18], PP1[18], PP2[18]);
  UBFA_18 U31 (W2[19], W6[18], PP3[18], PP4[18], PP5[18]);
  UBFA_18 U32 (W3[19], W7[18], PP6[18], PP7[18], PP8[18]);
  UBFA_18 U33 (W4[19], W8[18], PP9[18], PP10[18], PP11[18]);
  UBFA_19 U34 (W2[20], W5[19], PP0[19], PP1[19], PP2[19]);
  UBFA_19 U35 (W3[20], W6[19], PP3[19], PP4[19], PP5[19]);
  UBFA_19 U36 (W4[20], W7[19], PP6[19], PP7[19], PP8[19]);
  UBFA_19 U37 (W5[20], W8[19], PP9[19], PP10[19], PP11[19]);
  UBFA_20 U38 (W4[21], W6[20], PP0[20], PP1[20], PP2[20]);
  UBFA_20 U39 (W5[21], W7[20], PP3[20], PP4[20], PP5[20]);
  UBFA_20 U40 (W6[21], W8[20], PP6[20], PP7[20], PP8[20]);
  UBFA_21 U41 (W6[22], W7[21], PP0[21], PP1[21], PP2[21]);
  UBFA_21 U42 (W7[22], W8[21], PP3[21], PP4[21], PP5[21]);
  UBFA_22 U43 (W8[23], W8[22], PP0[22], PP1[22], PP2[22]);
  UBCON_8_0 U44 (W0[8:0], PP0[8:0]);
  UB1DCON_9 U45 (W0[9], PP2[9]);
  UB1DCON_10 U46 (W0[10], PP5[10]);
  UB1DCON_11 U47 (W0[11], PP8[11]);
  UB1DCON_12 U48 (W0[12], PP11[12]);
  UBCON_19_13 U49 (W0[19:13], PP12[19:13]);
  UB1DCON_20 U50 (W0[20], PP9[20]);
  UB1DCON_21 U51 (W0[21], PP6[21]);
  UB1DCON_22 U52 (W0[22], PP3[22]);
  UBCON_30_23 U53 (W0[30:23], PP0[30:23]);
  UBCON_8_1 U54 (W1[8:1], PP1[8:1]);
  UB1DCON_9 U55 (W1[9], PP3[9]);
  UB1DCON_10 U56 (W1[10], PP6[10]);
  UB1DCON_11 U57 (W1[11], PP9[11]);
  UB1DCON_12 U58 (W1[12], PP12[12]);
  UB1DCON_20 U59 (W1[20], PP10[20]);
  UB1DCON_21 U60 (W1[21], PP7[21]);
  UB1DCON_22 U61 (W1[22], PP4[22]);
  UBCON_29_23 U62 (W1[29:23], PP1[29:23]);
  UBCON_8_2 U63 (W2[8:2], PP2[8:2]);
  UB1DCON_9 U64 (W2[9], PP4[9]);
  UB1DCON_10 U65 (W2[10], PP7[10]);
  UB1DCON_11 U66 (W2[11], PP10[11]);
  UB1DCON_21 U67 (W2[21], PP8[21]);
  UB1DCON_22 U68 (W2[22], PP5[22]);
  UBCON_28_23 U69 (W2[28:23], PP2[28:23]);
  UBCON_8_3 U70 (W3[8:3], PP3[8:3]);
  UB1DCON_9 U71 (W3[9], PP5[9]);
  UB1DCON_10 U72 (W3[10], PP8[10]);
  UB1DCON_11 U73 (W3[11], PP11[11]);
  UB1DCON_21 U74 (W3[21], PP9[21]);
  UB1DCON_22 U75 (W3[22], PP6[22]);
  UBCON_27_23 U76 (W3[27:23], PP3[27:23]);
  UBCON_8_4 U77 (W4[8:4], PP4[8:4]);
  UB1DCON_9 U78 (W4[9], PP6[9]);
  UB1DCON_10 U79 (W4[10], PP9[10]);
  UB1DCON_22 U80 (W4[22], PP7[22]);
  UBCON_26_23 U81 (W4[26:23], PP4[26:23]);
  UBCON_8_5 U82 (W5[8:5], PP5[8:5]);
  UB1DCON_9 U83 (W5[9], PP7[9]);
  UB1DCON_10 U84 (W5[10], PP10[10]);
  UB1DCON_22 U85 (W5[22], PP8[22]);
  UBCON_25_23 U86 (W5[25:23], PP5[25:23]);
  UBCON_8_6 U87 (W6[8:6], PP6[8:6]);
  UB1DCON_9 U88 (W6[9], PP8[9]);
  UBCON_24_23 U89 (W6[24:23], PP6[24:23]);
  UBCON_8_7 U90 (W7[8:7], PP7[8:7]);
  UB1DCON_9 U91 (W7[9], PP9[9]);
  UB1DCON_23 U92 (W7[23], PP7[23]);
  UB1DCON_8 U93 (W8[8], PP8[8]);
  DADTR_30_0_29_1_2001 U94 (S1, S2, W0, W1, W2, W3, W4, W5, W6, W7, W8);
endmodule

module DADTR_30_0_29_1_2001 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8);
  output [30:0] S1;
  output [30:1] S2;
  input [30:0] PP0;
  input [29:1] PP1;
  input [28:2] PP2;
  input [27:3] PP3;
  input [26:4] PP4;
  input [25:5] PP5;
  input [24:6] PP6;
  input [23:7] PP7;
  input [23:8] PP8;
  wire [30:0] W0;
  wire [29:1] W1;
  wire [28:2] W2;
  wire [27:3] W3;
  wire [26:4] W4;
  wire [26:5] W5;
  UBHA_6 U0 (W3[7], W5[6], PP0[6], PP1[6]);
  UBFA_7 U1 (W1[8], W4[7], PP0[7], PP1[7], PP2[7]);
  UBHA_7 U2 (W2[8], W5[7], PP3[7], PP4[7]);
  UBFA_8 U3 (W0[9], W3[8], PP0[8], PP1[8], PP2[8]);
  UBFA_8 U4 (W1[9], W4[8], PP3[8], PP4[8], PP5[8]);
  UBHA_8 U5 (W2[9], W5[8], PP6[8], PP7[8]);
  UBFA_9 U6 (W0[10], W3[9], PP0[9], PP1[9], PP2[9]);
  UBFA_9 U7 (W1[10], W4[9], PP3[9], PP4[9], PP5[9]);
  UBFA_9 U8 (W2[10], W5[9], PP6[9], PP7[9], PP8[9]);
  UBFA_10 U9 (W0[11], W3[10], PP0[10], PP1[10], PP2[10]);
  UBFA_10 U10 (W1[11], W4[10], PP3[10], PP4[10], PP5[10]);
  UBFA_10 U11 (W2[11], W5[10], PP6[10], PP7[10], PP8[10]);
  UBFA_11 U12 (W0[12], W3[11], PP0[11], PP1[11], PP2[11]);
  UBFA_11 U13 (W1[12], W4[11], PP3[11], PP4[11], PP5[11]);
  UBFA_11 U14 (W2[12], W5[11], PP6[11], PP7[11], PP8[11]);
  UBFA_12 U15 (W0[13], W3[12], PP0[12], PP1[12], PP2[12]);
  UBFA_12 U16 (W1[13], W4[12], PP3[12], PP4[12], PP5[12]);
  UBFA_12 U17 (W2[13], W5[12], PP6[12], PP7[12], PP8[12]);
  UBFA_13 U18 (W0[14], W3[13], PP0[13], PP1[13], PP2[13]);
  UBFA_13 U19 (W1[14], W4[13], PP3[13], PP4[13], PP5[13]);
  UBFA_13 U20 (W2[14], W5[13], PP6[13], PP7[13], PP8[13]);
  UBFA_14 U21 (W0[15], W3[14], PP0[14], PP1[14], PP2[14]);
  UBFA_14 U22 (W1[15], W4[14], PP3[14], PP4[14], PP5[14]);
  UBFA_14 U23 (W2[15], W5[14], PP6[14], PP7[14], PP8[14]);
  UBFA_15 U24 (W0[16], W3[15], PP0[15], PP1[15], PP2[15]);
  UBFA_15 U25 (W1[16], W4[15], PP3[15], PP4[15], PP5[15]);
  UBFA_15 U26 (W2[16], W5[15], PP6[15], PP7[15], PP8[15]);
  UBFA_16 U27 (W0[17], W3[16], PP0[16], PP1[16], PP2[16]);
  UBFA_16 U28 (W1[17], W4[16], PP3[16], PP4[16], PP5[16]);
  UBFA_16 U29 (W2[17], W5[16], PP6[16], PP7[16], PP8[16]);
  UBFA_17 U30 (W0[18], W3[17], PP0[17], PP1[17], PP2[17]);
  UBFA_17 U31 (W1[18], W4[17], PP3[17], PP4[17], PP5[17]);
  UBFA_17 U32 (W2[18], W5[17], PP6[17], PP7[17], PP8[17]);
  UBFA_18 U33 (W0[19], W3[18], PP0[18], PP1[18], PP2[18]);
  UBFA_18 U34 (W1[19], W4[18], PP3[18], PP4[18], PP5[18]);
  UBFA_18 U35 (W2[19], W5[18], PP6[18], PP7[18], PP8[18]);
  UBFA_19 U36 (W0[20], W3[19], PP0[19], PP1[19], PP2[19]);
  UBFA_19 U37 (W1[20], W4[19], PP3[19], PP4[19], PP5[19]);
  UBFA_19 U38 (W2[20], W5[19], PP6[19], PP7[19], PP8[19]);
  UBFA_20 U39 (W0[21], W3[20], PP0[20], PP1[20], PP2[20]);
  UBFA_20 U40 (W1[21], W4[20], PP3[20], PP4[20], PP5[20]);
  UBFA_20 U41 (W2[21], W5[20], PP6[20], PP7[20], PP8[20]);
  UBFA_21 U42 (W0[22], W3[21], PP0[21], PP1[21], PP2[21]);
  UBFA_21 U43 (W1[22], W4[21], PP3[21], PP4[21], PP5[21]);
  UBFA_21 U44 (W2[22], W5[21], PP6[21], PP7[21], PP8[21]);
  UBFA_22 U45 (W0[23], W3[22], PP0[22], PP1[22], PP2[22]);
  UBFA_22 U46 (W1[23], W4[22], PP3[22], PP4[22], PP5[22]);
  UBFA_22 U47 (W2[23], W5[22], PP6[22], PP7[22], PP8[22]);
  UBFA_23 U48 (W1[24], W3[23], PP0[23], PP1[23], PP2[23]);
  UBFA_23 U49 (W2[24], W4[23], PP3[23], PP4[23], PP5[23]);
  UBFA_23 U50 (W3[24], W5[23], PP6[23], PP7[23], PP8[23]);
  UBFA_24 U51 (W3[25], W4[24], PP0[24], PP1[24], PP2[24]);
  UBFA_24 U52 (W4[25], W5[24], PP3[24], PP4[24], PP5[24]);
  UBFA_25 U53 (W5[26], W5[25], PP0[25], PP1[25], PP2[25]);
  UBCON_5_0 U54 (W0[5:0], PP0[5:0]);
  UB1DCON_6 U55 (W0[6], PP2[6]);
  UB1DCON_7 U56 (W0[7], PP5[7]);
  UB1DCON_8 U57 (W0[8], PP8[8]);
  UB1DCON_24 U58 (W0[24], PP6[24]);
  UB1DCON_25 U59 (W0[25], PP3[25]);
  UBCON_30_26 U60 (W0[30:26], PP0[30:26]);
  UBCON_5_1 U61 (W1[5:1], PP1[5:1]);
  UB1DCON_6 U62 (W1[6], PP3[6]);
  UB1DCON_7 U63 (W1[7], PP6[7]);
  UB1DCON_25 U64 (W1[25], PP4[25]);
  UBCON_29_26 U65 (W1[29:26], PP1[29:26]);
  UBCON_5_2 U66 (W2[5:2], PP2[5:2]);
  UB1DCON_6 U67 (W2[6], PP4[6]);
  UB1DCON_7 U68 (W2[7], PP7[7]);
  UB1DCON_25 U69 (W2[25], PP5[25]);
  UBCON_28_26 U70 (W2[28:26], PP2[28:26]);
  UBCON_5_3 U71 (W3[5:3], PP3[5:3]);
  UB1DCON_6 U72 (W3[6], PP5[6]);
  UBCON_27_26 U73 (W3[27:26], PP3[27:26]);
  UBCON_5_4 U74 (W4[5:4], PP4[5:4]);
  UB1DCON_6 U75 (W4[6], PP6[6]);
  UB1DCON_26 U76 (W4[26], PP4[26]);
  UB1DCON_5 U77 (W5[5], PP5[5]);
  DADTR_30_0_29_1_2002 U78 (S1, S2, W0, W1, W2, W3, W4, W5);
endmodule

module DADTR_30_0_29_1_2002 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5);
  output [30:0] S1;
  output [30:1] S2;
  input [30:0] PP0;
  input [29:1] PP1;
  input [28:2] PP2;
  input [27:3] PP3;
  input [26:4] PP4;
  input [26:5] PP5;
  wire [30:0] W0;
  wire [29:1] W1;
  wire [28:2] W2;
  wire [28:3] W3;
  UBHA_4 U0 (W1[5], W3[4], PP0[4], PP1[4]);
  UBFA_5 U1 (W0[6], W2[5], PP0[5], PP1[5], PP2[5]);
  UBHA_5 U2 (W1[6], W3[5], PP3[5], PP4[5]);
  UBFA_6 U3 (W0[7], W2[6], PP0[6], PP1[6], PP2[6]);
  UBFA_6 U4 (W1[7], W3[6], PP3[6], PP4[6], PP5[6]);
  UBFA_7 U5 (W0[8], W2[7], PP0[7], PP1[7], PP2[7]);
  UBFA_7 U6 (W1[8], W3[7], PP3[7], PP4[7], PP5[7]);
  UBFA_8 U7 (W0[9], W2[8], PP0[8], PP1[8], PP2[8]);
  UBFA_8 U8 (W1[9], W3[8], PP3[8], PP4[8], PP5[8]);
  UBFA_9 U9 (W0[10], W2[9], PP0[9], PP1[9], PP2[9]);
  UBFA_9 U10 (W1[10], W3[9], PP3[9], PP4[9], PP5[9]);
  UBFA_10 U11 (W0[11], W2[10], PP0[10], PP1[10], PP2[10]);
  UBFA_10 U12 (W1[11], W3[10], PP3[10], PP4[10], PP5[10]);
  UBFA_11 U13 (W0[12], W2[11], PP0[11], PP1[11], PP2[11]);
  UBFA_11 U14 (W1[12], W3[11], PP3[11], PP4[11], PP5[11]);
  UBFA_12 U15 (W0[13], W2[12], PP0[12], PP1[12], PP2[12]);
  UBFA_12 U16 (W1[13], W3[12], PP3[12], PP4[12], PP5[12]);
  UBFA_13 U17 (W0[14], W2[13], PP0[13], PP1[13], PP2[13]);
  UBFA_13 U18 (W1[14], W3[13], PP3[13], PP4[13], PP5[13]);
  UBFA_14 U19 (W0[15], W2[14], PP0[14], PP1[14], PP2[14]);
  UBFA_14 U20 (W1[15], W3[14], PP3[14], PP4[14], PP5[14]);
  UBFA_15 U21 (W0[16], W2[15], PP0[15], PP1[15], PP2[15]);
  UBFA_15 U22 (W1[16], W3[15], PP3[15], PP4[15], PP5[15]);
  UBFA_16 U23 (W0[17], W2[16], PP0[16], PP1[16], PP2[16]);
  UBFA_16 U24 (W1[17], W3[16], PP3[16], PP4[16], PP5[16]);
  UBFA_17 U25 (W0[18], W2[17], PP0[17], PP1[17], PP2[17]);
  UBFA_17 U26 (W1[18], W3[17], PP3[17], PP4[17], PP5[17]);
  UBFA_18 U27 (W0[19], W2[18], PP0[18], PP1[18], PP2[18]);
  UBFA_18 U28 (W1[19], W3[18], PP3[18], PP4[18], PP5[18]);
  UBFA_19 U29 (W0[20], W2[19], PP0[19], PP1[19], PP2[19]);
  UBFA_19 U30 (W1[20], W3[19], PP3[19], PP4[19], PP5[19]);
  UBFA_20 U31 (W0[21], W2[20], PP0[20], PP1[20], PP2[20]);
  UBFA_20 U32 (W1[21], W3[20], PP3[20], PP4[20], PP5[20]);
  UBFA_21 U33 (W0[22], W2[21], PP0[21], PP1[21], PP2[21]);
  UBFA_21 U34 (W1[22], W3[21], PP3[21], PP4[21], PP5[21]);
  UBFA_22 U35 (W0[23], W2[22], PP0[22], PP1[22], PP2[22]);
  UBFA_22 U36 (W1[23], W3[22], PP3[22], PP4[22], PP5[22]);
  UBFA_23 U37 (W0[24], W2[23], PP0[23], PP1[23], PP2[23]);
  UBFA_23 U38 (W1[24], W3[23], PP3[23], PP4[23], PP5[23]);
  UBFA_24 U39 (W0[25], W2[24], PP0[24], PP1[24], PP2[24]);
  UBFA_24 U40 (W1[25], W3[24], PP3[24], PP4[24], PP5[24]);
  UBFA_25 U41 (W0[26], W2[25], PP0[25], PP1[25], PP2[25]);
  UBFA_25 U42 (W1[26], W3[25], PP3[25], PP4[25], PP5[25]);
  UBFA_26 U43 (W1[27], W2[26], PP0[26], PP1[26], PP2[26]);
  UBFA_26 U44 (W2[27], W3[26], PP3[26], PP4[26], PP5[26]);
  UBFA_27 U45 (W3[28], W3[27], PP0[27], PP1[27], PP2[27]);
  UBCON_3_0 U46 (W0[3:0], PP0[3:0]);
  UB1DCON_4 U47 (W0[4], PP2[4]);
  UB1DCON_5 U48 (W0[5], PP5[5]);
  UB1DCON_27 U49 (W0[27], PP3[27]);
  UBCON_30_28 U50 (W0[30:28], PP0[30:28]);
  UBCON_3_1 U51 (W1[3:1], PP1[3:1]);
  UB1DCON_4 U52 (W1[4], PP3[4]);
  UBCON_29_28 U53 (W1[29:28], PP1[29:28]);
  UBCON_3_2 U54 (W2[3:2], PP2[3:2]);
  UB1DCON_4 U55 (W2[4], PP4[4]);
  UB1DCON_28 U56 (W2[28], PP2[28]);
  UB1DCON_3 U57 (W3[3], PP3[3]);
  DADTR_30_0_29_1_2003 U58 (S1, S2, W0, W1, W2, W3);
endmodule

module DADTR_30_0_29_1_2003 (S1, S2, PP0, PP1, PP2, PP3);
  output [30:0] S1;
  output [30:1] S2;
  input [30:0] PP0;
  input [29:1] PP1;
  input [28:2] PP2;
  input [28:3] PP3;
  wire [30:0] W0;
  wire [29:1] W1;
  wire [29:2] W2;
  UBHA_3 U0 (W1[4], W2[3], PP0[3], PP1[3]);
  UBFA_4 U1 (W1[5], W2[4], PP0[4], PP1[4], PP2[4]);
  UBFA_5 U2 (W1[6], W2[5], PP0[5], PP1[5], PP2[5]);
  UBFA_6 U3 (W1[7], W2[6], PP0[6], PP1[6], PP2[6]);
  UBFA_7 U4 (W1[8], W2[7], PP0[7], PP1[7], PP2[7]);
  UBFA_8 U5 (W1[9], W2[8], PP0[8], PP1[8], PP2[8]);
  UBFA_9 U6 (W1[10], W2[9], PP0[9], PP1[9], PP2[9]);
  UBFA_10 U7 (W1[11], W2[10], PP0[10], PP1[10], PP2[10]);
  UBFA_11 U8 (W1[12], W2[11], PP0[11], PP1[11], PP2[11]);
  UBFA_12 U9 (W1[13], W2[12], PP0[12], PP1[12], PP2[12]);
  UBFA_13 U10 (W1[14], W2[13], PP0[13], PP1[13], PP2[13]);
  UBFA_14 U11 (W1[15], W2[14], PP0[14], PP1[14], PP2[14]);
  UBFA_15 U12 (W1[16], W2[15], PP0[15], PP1[15], PP2[15]);
  UBFA_16 U13 (W1[17], W2[16], PP0[16], PP1[16], PP2[16]);
  UBFA_17 U14 (W1[18], W2[17], PP0[17], PP1[17], PP2[17]);
  UBFA_18 U15 (W1[19], W2[18], PP0[18], PP1[18], PP2[18]);
  UBFA_19 U16 (W1[20], W2[19], PP0[19], PP1[19], PP2[19]);
  UBFA_20 U17 (W1[21], W2[20], PP0[20], PP1[20], PP2[20]);
  UBFA_21 U18 (W1[22], W2[21], PP0[21], PP1[21], PP2[21]);
  UBFA_22 U19 (W1[23], W2[22], PP0[22], PP1[22], PP2[22]);
  UBFA_23 U20 (W1[24], W2[23], PP0[23], PP1[23], PP2[23]);
  UBFA_24 U21 (W1[25], W2[24], PP0[24], PP1[24], PP2[24]);
  UBFA_25 U22 (W1[26], W2[25], PP0[25], PP1[25], PP2[25]);
  UBFA_26 U23 (W1[27], W2[26], PP0[26], PP1[26], PP2[26]);
  UBFA_27 U24 (W1[28], W2[27], PP0[27], PP1[27], PP2[27]);
  UBFA_28 U25 (W2[29], W2[28], PP0[28], PP1[28], PP2[28]);
  UBCON_2_0 U26 (W0[2:0], PP0[2:0]);
  UB1DCON_3 U27 (W0[3], PP2[3]);
  UBCON_28_4 U28 (W0[28:4], PP3[28:4]);
  UBCON_30_29 U29 (W0[30:29], PP0[30:29]);
  UBCON_2_1 U30 (W1[2:1], PP1[2:1]);
  UB1DCON_3 U31 (W1[3], PP3[3]);
  UB1DCON_29 U32 (W1[29], PP1[29]);
  UB1DCON_2 U33 (W2[2], PP2[2]);
  DADTR_30_0_29_1_2004 U34 (S1, S2, W0, W1, W2);
endmodule

module DADTR_30_0_29_1_2004 (S1, S2, PP0, PP1, PP2);
  output [30:0] S1;
  output [30:1] S2;
  input [30:0] PP0;
  input [29:1] PP1;
  input [29:2] PP2;
  wire [30:0] W0;
  wire [30:1] W1;
  UBHA_2 U0 (W0[3], W1[2], PP0[2], PP1[2]);
  UBFA_3 U1 (W0[4], W1[3], PP0[3], PP1[3], PP2[3]);
  UBFA_4 U2 (W0[5], W1[4], PP0[4], PP1[4], PP2[4]);
  UBFA_5 U3 (W0[6], W1[5], PP0[5], PP1[5], PP2[5]);
  UBFA_6 U4 (W0[7], W1[6], PP0[6], PP1[6], PP2[6]);
  UBFA_7 U5 (W0[8], W1[7], PP0[7], PP1[7], PP2[7]);
  UBFA_8 U6 (W0[9], W1[8], PP0[8], PP1[8], PP2[8]);
  UBFA_9 U7 (W0[10], W1[9], PP0[9], PP1[9], PP2[9]);
  UBFA_10 U8 (W0[11], W1[10], PP0[10], PP1[10], PP2[10]);
  UBFA_11 U9 (W0[12], W1[11], PP0[11], PP1[11], PP2[11]);
  UBFA_12 U10 (W0[13], W1[12], PP0[12], PP1[12], PP2[12]);
  UBFA_13 U11 (W0[14], W1[13], PP0[13], PP1[13], PP2[13]);
  UBFA_14 U12 (W0[15], W1[14], PP0[14], PP1[14], PP2[14]);
  UBFA_15 U13 (W0[16], W1[15], PP0[15], PP1[15], PP2[15]);
  UBFA_16 U14 (W0[17], W1[16], PP0[16], PP1[16], PP2[16]);
  UBFA_17 U15 (W0[18], W1[17], PP0[17], PP1[17], PP2[17]);
  UBFA_18 U16 (W0[19], W1[18], PP0[18], PP1[18], PP2[18]);
  UBFA_19 U17 (W0[20], W1[19], PP0[19], PP1[19], PP2[19]);
  UBFA_20 U18 (W0[21], W1[20], PP0[20], PP1[20], PP2[20]);
  UBFA_21 U19 (W0[22], W1[21], PP0[21], PP1[21], PP2[21]);
  UBFA_22 U20 (W0[23], W1[22], PP0[22], PP1[22], PP2[22]);
  UBFA_23 U21 (W0[24], W1[23], PP0[23], PP1[23], PP2[23]);
  UBFA_24 U22 (W0[25], W1[24], PP0[24], PP1[24], PP2[24]);
  UBFA_25 U23 (W0[26], W1[25], PP0[25], PP1[25], PP2[25]);
  UBFA_26 U24 (W0[27], W1[26], PP0[26], PP1[26], PP2[26]);
  UBFA_27 U25 (W0[28], W1[27], PP0[27], PP1[27], PP2[27]);
  UBFA_28 U26 (W0[29], W1[28], PP0[28], PP1[28], PP2[28]);
  UBFA_29 U27 (W1[30], W1[29], PP0[29], PP1[29], PP2[29]);
  UBCON_1_0 U28 (W0[1:0], PP0[1:0]);
  UB1DCON_2 U29 (W0[2], PP2[2]);
  UB1DCON_30 U30 (W0[30], PP0[30]);
  UB1DCON_1 U31 (W1[1], PP1[1]);
  DADTR_30_0_30_1 U32 (S1, S2, W0, W1);
endmodule

module DADTR_30_0_30_1 (S1, S2, PP0, PP1);
  output [30:0] S1;
  output [30:1] S2;
  input [30:0] PP0;
  input [30:1] PP1;
  UBCON_30_0 U0 (S1, PP0);
  UBCON_30_1 U1 (S2, PP1);
endmodule

module MultUB_STD_DAD_KS000 (P, IN1, IN2);
  output [31:0] P;
  input [15:0] IN1;
  input [15:0] IN2;
  wire [15:0] PP0;
  wire [16:1] PP1;
  wire [25:10] PP10;
  wire [26:11] PP11;
  wire [27:12] PP12;
  wire [28:13] PP13;
  wire [29:14] PP14;
  wire [30:15] PP15;
  wire [17:2] PP2;
  wire [18:3] PP3;
  wire [19:4] PP4;
  wire [20:5] PP5;
  wire [21:6] PP6;
  wire [22:7] PP7;
  wire [23:8] PP8;
  wire [24:9] PP9;
  wire [30:0] S1;
  wire [30:1] S2;
  UBPPG_15_0_15_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, IN1, IN2);
  DADTR_15_0_16_1_1000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15);
  UBKSA_30_0_30_1 U2 (P, S1, S2);
endmodule

module UBCON_12_0 (O, I);
  output [12:0] O;
  input [12:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
endmodule

module UBCON_12_1 (O, I);
  output [12:1] O;
  input [12:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
  UB1DCON_6 U5 (O[6], I[6]);
  UB1DCON_7 U6 (O[7], I[7]);
  UB1DCON_8 U7 (O[8], I[8]);
  UB1DCON_9 U8 (O[9], I[9]);
  UB1DCON_10 U9 (O[10], I[10]);
  UB1DCON_11 U10 (O[11], I[11]);
  UB1DCON_12 U11 (O[12], I[12]);
endmodule

module UBCON_12_10 (O, I);
  output [12:10] O;
  input [12:10] I;
  UB1DCON_10 U0 (O[10], I[10]);
  UB1DCON_11 U1 (O[11], I[11]);
  UB1DCON_12 U2 (O[12], I[12]);
endmodule

module UBCON_12_11 (O, I);
  output [12:11] O;
  input [12:11] I;
  UB1DCON_11 U0 (O[11], I[11]);
  UB1DCON_12 U1 (O[12], I[12]);
endmodule

module UBCON_12_2 (O, I);
  output [12:2] O;
  input [12:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
  UB1DCON_6 U4 (O[6], I[6]);
  UB1DCON_7 U5 (O[7], I[7]);
  UB1DCON_8 U6 (O[8], I[8]);
  UB1DCON_9 U7 (O[9], I[9]);
  UB1DCON_10 U8 (O[10], I[10]);
  UB1DCON_11 U9 (O[11], I[11]);
  UB1DCON_12 U10 (O[12], I[12]);
endmodule

module UBCON_12_3 (O, I);
  output [12:3] O;
  input [12:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
  UB1DCON_6 U3 (O[6], I[6]);
  UB1DCON_7 U4 (O[7], I[7]);
  UB1DCON_8 U5 (O[8], I[8]);
  UB1DCON_9 U6 (O[9], I[9]);
  UB1DCON_10 U7 (O[10], I[10]);
  UB1DCON_11 U8 (O[11], I[11]);
  UB1DCON_12 U9 (O[12], I[12]);
endmodule

module UBCON_12_4 (O, I);
  output [12:4] O;
  input [12:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
  UB1DCON_11 U7 (O[11], I[11]);
  UB1DCON_12 U8 (O[12], I[12]);
endmodule

module UBCON_12_5 (O, I);
  output [12:5] O;
  input [12:5] I;
  UB1DCON_5 U0 (O[5], I[5]);
  UB1DCON_6 U1 (O[6], I[6]);
  UB1DCON_7 U2 (O[7], I[7]);
  UB1DCON_8 U3 (O[8], I[8]);
  UB1DCON_9 U4 (O[9], I[9]);
  UB1DCON_10 U5 (O[10], I[10]);
  UB1DCON_11 U6 (O[11], I[11]);
  UB1DCON_12 U7 (O[12], I[12]);
endmodule

module UBCON_12_6 (O, I);
  output [12:6] O;
  input [12:6] I;
  UB1DCON_6 U0 (O[6], I[6]);
  UB1DCON_7 U1 (O[7], I[7]);
  UB1DCON_8 U2 (O[8], I[8]);
  UB1DCON_9 U3 (O[9], I[9]);
  UB1DCON_10 U4 (O[10], I[10]);
  UB1DCON_11 U5 (O[11], I[11]);
  UB1DCON_12 U6 (O[12], I[12]);
endmodule

module UBCON_12_7 (O, I);
  output [12:7] O;
  input [12:7] I;
  UB1DCON_7 U0 (O[7], I[7]);
  UB1DCON_8 U1 (O[8], I[8]);
  UB1DCON_9 U2 (O[9], I[9]);
  UB1DCON_10 U3 (O[10], I[10]);
  UB1DCON_11 U4 (O[11], I[11]);
  UB1DCON_12 U5 (O[12], I[12]);
endmodule

module UBCON_12_8 (O, I);
  output [12:8] O;
  input [12:8] I;
  UB1DCON_8 U0 (O[8], I[8]);
  UB1DCON_9 U1 (O[9], I[9]);
  UB1DCON_10 U2 (O[10], I[10]);
  UB1DCON_11 U3 (O[11], I[11]);
  UB1DCON_12 U4 (O[12], I[12]);
endmodule

module UBCON_12_9 (O, I);
  output [12:9] O;
  input [12:9] I;
  UB1DCON_9 U0 (O[9], I[9]);
  UB1DCON_10 U1 (O[10], I[10]);
  UB1DCON_11 U2 (O[11], I[11]);
  UB1DCON_12 U3 (O[12], I[12]);
endmodule

module UBCON_19_13 (O, I);
  output [19:13] O;
  input [19:13] I;
  UB1DCON_13 U0 (O[13], I[13]);
  UB1DCON_14 U1 (O[14], I[14]);
  UB1DCON_15 U2 (O[15], I[15]);
  UB1DCON_16 U3 (O[16], I[16]);
  UB1DCON_17 U4 (O[17], I[17]);
  UB1DCON_18 U5 (O[18], I[18]);
  UB1DCON_19 U6 (O[19], I[19]);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_24_23 (O, I);
  output [24:23] O;
  input [24:23] I;
  UB1DCON_23 U0 (O[23], I[23]);
  UB1DCON_24 U1 (O[24], I[24]);
endmodule

module UBCON_25_23 (O, I);
  output [25:23] O;
  input [25:23] I;
  UB1DCON_23 U0 (O[23], I[23]);
  UB1DCON_24 U1 (O[24], I[24]);
  UB1DCON_25 U2 (O[25], I[25]);
endmodule

module UBCON_26_23 (O, I);
  output [26:23] O;
  input [26:23] I;
  UB1DCON_23 U0 (O[23], I[23]);
  UB1DCON_24 U1 (O[24], I[24]);
  UB1DCON_25 U2 (O[25], I[25]);
  UB1DCON_26 U3 (O[26], I[26]);
endmodule

module UBCON_27_23 (O, I);
  output [27:23] O;
  input [27:23] I;
  UB1DCON_23 U0 (O[23], I[23]);
  UB1DCON_24 U1 (O[24], I[24]);
  UB1DCON_25 U2 (O[25], I[25]);
  UB1DCON_26 U3 (O[26], I[26]);
  UB1DCON_27 U4 (O[27], I[27]);
endmodule

module UBCON_27_26 (O, I);
  output [27:26] O;
  input [27:26] I;
  UB1DCON_26 U0 (O[26], I[26]);
  UB1DCON_27 U1 (O[27], I[27]);
endmodule

module UBCON_28_23 (O, I);
  output [28:23] O;
  input [28:23] I;
  UB1DCON_23 U0 (O[23], I[23]);
  UB1DCON_24 U1 (O[24], I[24]);
  UB1DCON_25 U2 (O[25], I[25]);
  UB1DCON_26 U3 (O[26], I[26]);
  UB1DCON_27 U4 (O[27], I[27]);
  UB1DCON_28 U5 (O[28], I[28]);
endmodule

module UBCON_28_26 (O, I);
  output [28:26] O;
  input [28:26] I;
  UB1DCON_26 U0 (O[26], I[26]);
  UB1DCON_27 U1 (O[27], I[27]);
  UB1DCON_28 U2 (O[28], I[28]);
endmodule

module UBCON_28_4 (O, I);
  output [28:4] O;
  input [28:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
  UB1DCON_9 U5 (O[9], I[9]);
  UB1DCON_10 U6 (O[10], I[10]);
  UB1DCON_11 U7 (O[11], I[11]);
  UB1DCON_12 U8 (O[12], I[12]);
  UB1DCON_13 U9 (O[13], I[13]);
  UB1DCON_14 U10 (O[14], I[14]);
  UB1DCON_15 U11 (O[15], I[15]);
  UB1DCON_16 U12 (O[16], I[16]);
  UB1DCON_17 U13 (O[17], I[17]);
  UB1DCON_18 U14 (O[18], I[18]);
  UB1DCON_19 U15 (O[19], I[19]);
  UB1DCON_20 U16 (O[20], I[20]);
  UB1DCON_21 U17 (O[21], I[21]);
  UB1DCON_22 U18 (O[22], I[22]);
  UB1DCON_23 U19 (O[23], I[23]);
  UB1DCON_24 U20 (O[24], I[24]);
  UB1DCON_25 U21 (O[25], I[25]);
  UB1DCON_26 U22 (O[26], I[26]);
  UB1DCON_27 U23 (O[27], I[27]);
  UB1DCON_28 U24 (O[28], I[28]);
endmodule

module UBCON_29_23 (O, I);
  output [29:23] O;
  input [29:23] I;
  UB1DCON_23 U0 (O[23], I[23]);
  UB1DCON_24 U1 (O[24], I[24]);
  UB1DCON_25 U2 (O[25], I[25]);
  UB1DCON_26 U3 (O[26], I[26]);
  UB1DCON_27 U4 (O[27], I[27]);
  UB1DCON_28 U5 (O[28], I[28]);
  UB1DCON_29 U6 (O[29], I[29]);
endmodule

module UBCON_29_26 (O, I);
  output [29:26] O;
  input [29:26] I;
  UB1DCON_26 U0 (O[26], I[26]);
  UB1DCON_27 U1 (O[27], I[27]);
  UB1DCON_28 U2 (O[28], I[28]);
  UB1DCON_29 U3 (O[29], I[29]);
endmodule

module UBCON_29_28 (O, I);
  output [29:28] O;
  input [29:28] I;
  UB1DCON_28 U0 (O[28], I[28]);
  UB1DCON_29 U1 (O[29], I[29]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBCON_2_1 (O, I);
  output [2:1] O;
  input [2:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
endmodule

module UBCON_30_0 (O, I);
  output [30:0] O;
  input [30:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
  UB1DCON_13 U13 (O[13], I[13]);
  UB1DCON_14 U14 (O[14], I[14]);
  UB1DCON_15 U15 (O[15], I[15]);
  UB1DCON_16 U16 (O[16], I[16]);
  UB1DCON_17 U17 (O[17], I[17]);
  UB1DCON_18 U18 (O[18], I[18]);
  UB1DCON_19 U19 (O[19], I[19]);
  UB1DCON_20 U20 (O[20], I[20]);
  UB1DCON_21 U21 (O[21], I[21]);
  UB1DCON_22 U22 (O[22], I[22]);
  UB1DCON_23 U23 (O[23], I[23]);
  UB1DCON_24 U24 (O[24], I[24]);
  UB1DCON_25 U25 (O[25], I[25]);
  UB1DCON_26 U26 (O[26], I[26]);
  UB1DCON_27 U27 (O[27], I[27]);
  UB1DCON_28 U28 (O[28], I[28]);
  UB1DCON_29 U29 (O[29], I[29]);
  UB1DCON_30 U30 (O[30], I[30]);
endmodule

module UBCON_30_1 (O, I);
  output [30:1] O;
  input [30:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
  UB1DCON_6 U5 (O[6], I[6]);
  UB1DCON_7 U6 (O[7], I[7]);
  UB1DCON_8 U7 (O[8], I[8]);
  UB1DCON_9 U8 (O[9], I[9]);
  UB1DCON_10 U9 (O[10], I[10]);
  UB1DCON_11 U10 (O[11], I[11]);
  UB1DCON_12 U11 (O[12], I[12]);
  UB1DCON_13 U12 (O[13], I[13]);
  UB1DCON_14 U13 (O[14], I[14]);
  UB1DCON_15 U14 (O[15], I[15]);
  UB1DCON_16 U15 (O[16], I[16]);
  UB1DCON_17 U16 (O[17], I[17]);
  UB1DCON_18 U17 (O[18], I[18]);
  UB1DCON_19 U18 (O[19], I[19]);
  UB1DCON_20 U19 (O[20], I[20]);
  UB1DCON_21 U20 (O[21], I[21]);
  UB1DCON_22 U21 (O[22], I[22]);
  UB1DCON_23 U22 (O[23], I[23]);
  UB1DCON_24 U23 (O[24], I[24]);
  UB1DCON_25 U24 (O[25], I[25]);
  UB1DCON_26 U25 (O[26], I[26]);
  UB1DCON_27 U26 (O[27], I[27]);
  UB1DCON_28 U27 (O[28], I[28]);
  UB1DCON_29 U28 (O[29], I[29]);
  UB1DCON_30 U29 (O[30], I[30]);
endmodule

module UBCON_30_23 (O, I);
  output [30:23] O;
  input [30:23] I;
  UB1DCON_23 U0 (O[23], I[23]);
  UB1DCON_24 U1 (O[24], I[24]);
  UB1DCON_25 U2 (O[25], I[25]);
  UB1DCON_26 U3 (O[26], I[26]);
  UB1DCON_27 U4 (O[27], I[27]);
  UB1DCON_28 U5 (O[28], I[28]);
  UB1DCON_29 U6 (O[29], I[29]);
  UB1DCON_30 U7 (O[30], I[30]);
endmodule

module UBCON_30_26 (O, I);
  output [30:26] O;
  input [30:26] I;
  UB1DCON_26 U0 (O[26], I[26]);
  UB1DCON_27 U1 (O[27], I[27]);
  UB1DCON_28 U2 (O[28], I[28]);
  UB1DCON_29 U3 (O[29], I[29]);
  UB1DCON_30 U4 (O[30], I[30]);
endmodule

module UBCON_30_28 (O, I);
  output [30:28] O;
  input [30:28] I;
  UB1DCON_28 U0 (O[28], I[28]);
  UB1DCON_29 U1 (O[29], I[29]);
  UB1DCON_30 U2 (O[30], I[30]);
endmodule

module UBCON_30_29 (O, I);
  output [30:29] O;
  input [30:29] I;
  UB1DCON_29 U0 (O[29], I[29]);
  UB1DCON_30 U1 (O[30], I[30]);
endmodule

module UBCON_3_0 (O, I);
  output [3:0] O;
  input [3:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
endmodule

module UBCON_3_1 (O, I);
  output [3:1] O;
  input [3:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
endmodule

module UBCON_3_2 (O, I);
  output [3:2] O;
  input [3:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
endmodule

module UBCON_5_0 (O, I);
  output [5:0] O;
  input [5:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
endmodule

module UBCON_5_1 (O, I);
  output [5:1] O;
  input [5:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
endmodule

module UBCON_5_2 (O, I);
  output [5:2] O;
  input [5:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
endmodule

module UBCON_5_3 (O, I);
  output [5:3] O;
  input [5:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
endmodule

module UBCON_5_4 (O, I);
  output [5:4] O;
  input [5:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
endmodule

module UBCON_8_0 (O, I);
  output [8:0] O;
  input [8:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
endmodule

module UBCON_8_1 (O, I);
  output [8:1] O;
  input [8:1] I;
  UB1DCON_1 U0 (O[1], I[1]);
  UB1DCON_2 U1 (O[2], I[2]);
  UB1DCON_3 U2 (O[3], I[3]);
  UB1DCON_4 U3 (O[4], I[4]);
  UB1DCON_5 U4 (O[5], I[5]);
  UB1DCON_6 U5 (O[6], I[6]);
  UB1DCON_7 U6 (O[7], I[7]);
  UB1DCON_8 U7 (O[8], I[8]);
endmodule

module UBCON_8_2 (O, I);
  output [8:2] O;
  input [8:2] I;
  UB1DCON_2 U0 (O[2], I[2]);
  UB1DCON_3 U1 (O[3], I[3]);
  UB1DCON_4 U2 (O[4], I[4]);
  UB1DCON_5 U3 (O[5], I[5]);
  UB1DCON_6 U4 (O[6], I[6]);
  UB1DCON_7 U5 (O[7], I[7]);
  UB1DCON_8 U6 (O[8], I[8]);
endmodule

module UBCON_8_3 (O, I);
  output [8:3] O;
  input [8:3] I;
  UB1DCON_3 U0 (O[3], I[3]);
  UB1DCON_4 U1 (O[4], I[4]);
  UB1DCON_5 U2 (O[5], I[5]);
  UB1DCON_6 U3 (O[6], I[6]);
  UB1DCON_7 U4 (O[7], I[7]);
  UB1DCON_8 U5 (O[8], I[8]);
endmodule

module UBCON_8_4 (O, I);
  output [8:4] O;
  input [8:4] I;
  UB1DCON_4 U0 (O[4], I[4]);
  UB1DCON_5 U1 (O[5], I[5]);
  UB1DCON_6 U2 (O[6], I[6]);
  UB1DCON_7 U3 (O[7], I[7]);
  UB1DCON_8 U4 (O[8], I[8]);
endmodule

module UBCON_8_5 (O, I);
  output [8:5] O;
  input [8:5] I;
  UB1DCON_5 U0 (O[5], I[5]);
  UB1DCON_6 U1 (O[6], I[6]);
  UB1DCON_7 U2 (O[7], I[7]);
  UB1DCON_8 U3 (O[8], I[8]);
endmodule

module UBCON_8_6 (O, I);
  output [8:6] O;
  input [8:6] I;
  UB1DCON_6 U0 (O[6], I[6]);
  UB1DCON_7 U1 (O[7], I[7]);
  UB1DCON_8 U2 (O[8], I[8]);
endmodule

module UBCON_8_7 (O, I);
  output [8:7] O;
  input [8:7] I;
  UB1DCON_7 U0 (O[7], I[7]);
  UB1DCON_8 U1 (O[8], I[8]);
endmodule

module UBKSA_30_0_30_1 (S, X, Y);
  output [31:0] S;
  input [30:0] X;
  input [30:1] Y;
  UBPureKSA_30_1 U0 (S[31:1], X[30:1], Y[30:1]);
  UB1DCON_0 U1 (S[0], X[0]);
endmodule

module UBPPG_15_0_15_0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, IN1, IN2);
  output [15:0] PP0;
  output [16:1] PP1;
  output [25:10] PP10;
  output [26:11] PP11;
  output [27:12] PP12;
  output [28:13] PP13;
  output [29:14] PP14;
  output [30:15] PP15;
  output [17:2] PP2;
  output [18:3] PP3;
  output [19:4] PP4;
  output [20:5] PP5;
  output [21:6] PP6;
  output [22:7] PP7;
  output [23:8] PP8;
  output [24:9] PP9;
  input [15:0] IN1;
  input [15:0] IN2;
  UBVPPG_15_0_0 U0 (PP0, IN1, IN2[0]);
  UBVPPG_15_0_1 U1 (PP1, IN1, IN2[1]);
  UBVPPG_15_0_2 U2 (PP2, IN1, IN2[2]);
  UBVPPG_15_0_3 U3 (PP3, IN1, IN2[3]);
  UBVPPG_15_0_4 U4 (PP4, IN1, IN2[4]);
  UBVPPG_15_0_5 U5 (PP5, IN1, IN2[5]);
  UBVPPG_15_0_6 U6 (PP6, IN1, IN2[6]);
  UBVPPG_15_0_7 U7 (PP7, IN1, IN2[7]);
  UBVPPG_15_0_8 U8 (PP8, IN1, IN2[8]);
  UBVPPG_15_0_9 U9 (PP9, IN1, IN2[9]);
  UBVPPG_15_0_10 U10 (PP10, IN1, IN2[10]);
  UBVPPG_15_0_11 U11 (PP11, IN1, IN2[11]);
  UBVPPG_15_0_12 U12 (PP12, IN1, IN2[12]);
  UBVPPG_15_0_13 U13 (PP13, IN1, IN2[13]);
  UBVPPG_15_0_14 U14 (PP14, IN1, IN2[14]);
  UBVPPG_15_0_15 U15 (PP15, IN1, IN2[15]);
endmodule

module UBPureKSA_30_1 (S, X, Y);
  output [31:1] S;
  input [30:1] X;
  input [30:1] Y;
  wire C;
  UBPriKSA_30_1 U0 (S, X, Y, C);
  UBZero_1_1 U1 (C);
endmodule

module UBVPPG_15_0_0 (O, IN1, IN2);
  output [15:0] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_0 U0 (O[0], IN1[0], IN2);
  UB1BPPG_1_0 U1 (O[1], IN1[1], IN2);
  UB1BPPG_2_0 U2 (O[2], IN1[2], IN2);
  UB1BPPG_3_0 U3 (O[3], IN1[3], IN2);
  UB1BPPG_4_0 U4 (O[4], IN1[4], IN2);
  UB1BPPG_5_0 U5 (O[5], IN1[5], IN2);
  UB1BPPG_6_0 U6 (O[6], IN1[6], IN2);
  UB1BPPG_7_0 U7 (O[7], IN1[7], IN2);
  UB1BPPG_8_0 U8 (O[8], IN1[8], IN2);
  UB1BPPG_9_0 U9 (O[9], IN1[9], IN2);
  UB1BPPG_10_0 U10 (O[10], IN1[10], IN2);
  UB1BPPG_11_0 U11 (O[11], IN1[11], IN2);
  UB1BPPG_12_0 U12 (O[12], IN1[12], IN2);
  UB1BPPG_13_0 U13 (O[13], IN1[13], IN2);
  UB1BPPG_14_0 U14 (O[14], IN1[14], IN2);
  UB1BPPG_15_0 U15 (O[15], IN1[15], IN2);
endmodule

module UBVPPG_15_0_1 (O, IN1, IN2);
  output [16:1] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_1 U0 (O[1], IN1[0], IN2);
  UB1BPPG_1_1 U1 (O[2], IN1[1], IN2);
  UB1BPPG_2_1 U2 (O[3], IN1[2], IN2);
  UB1BPPG_3_1 U3 (O[4], IN1[3], IN2);
  UB1BPPG_4_1 U4 (O[5], IN1[4], IN2);
  UB1BPPG_5_1 U5 (O[6], IN1[5], IN2);
  UB1BPPG_6_1 U6 (O[7], IN1[6], IN2);
  UB1BPPG_7_1 U7 (O[8], IN1[7], IN2);
  UB1BPPG_8_1 U8 (O[9], IN1[8], IN2);
  UB1BPPG_9_1 U9 (O[10], IN1[9], IN2);
  UB1BPPG_10_1 U10 (O[11], IN1[10], IN2);
  UB1BPPG_11_1 U11 (O[12], IN1[11], IN2);
  UB1BPPG_12_1 U12 (O[13], IN1[12], IN2);
  UB1BPPG_13_1 U13 (O[14], IN1[13], IN2);
  UB1BPPG_14_1 U14 (O[15], IN1[14], IN2);
  UB1BPPG_15_1 U15 (O[16], IN1[15], IN2);
endmodule

module UBVPPG_15_0_10 (O, IN1, IN2);
  output [25:10] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_10 U0 (O[10], IN1[0], IN2);
  UB1BPPG_1_10 U1 (O[11], IN1[1], IN2);
  UB1BPPG_2_10 U2 (O[12], IN1[2], IN2);
  UB1BPPG_3_10 U3 (O[13], IN1[3], IN2);
  UB1BPPG_4_10 U4 (O[14], IN1[4], IN2);
  UB1BPPG_5_10 U5 (O[15], IN1[5], IN2);
  UB1BPPG_6_10 U6 (O[16], IN1[6], IN2);
  UB1BPPG_7_10 U7 (O[17], IN1[7], IN2);
  UB1BPPG_8_10 U8 (O[18], IN1[8], IN2);
  UB1BPPG_9_10 U9 (O[19], IN1[9], IN2);
  UB1BPPG_10_10 U10 (O[20], IN1[10], IN2);
  UB1BPPG_11_10 U11 (O[21], IN1[11], IN2);
  UB1BPPG_12_10 U12 (O[22], IN1[12], IN2);
  UB1BPPG_13_10 U13 (O[23], IN1[13], IN2);
  UB1BPPG_14_10 U14 (O[24], IN1[14], IN2);
  UB1BPPG_15_10 U15 (O[25], IN1[15], IN2);
endmodule

module UBVPPG_15_0_11 (O, IN1, IN2);
  output [26:11] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_11 U0 (O[11], IN1[0], IN2);
  UB1BPPG_1_11 U1 (O[12], IN1[1], IN2);
  UB1BPPG_2_11 U2 (O[13], IN1[2], IN2);
  UB1BPPG_3_11 U3 (O[14], IN1[3], IN2);
  UB1BPPG_4_11 U4 (O[15], IN1[4], IN2);
  UB1BPPG_5_11 U5 (O[16], IN1[5], IN2);
  UB1BPPG_6_11 U6 (O[17], IN1[6], IN2);
  UB1BPPG_7_11 U7 (O[18], IN1[7], IN2);
  UB1BPPG_8_11 U8 (O[19], IN1[8], IN2);
  UB1BPPG_9_11 U9 (O[20], IN1[9], IN2);
  UB1BPPG_10_11 U10 (O[21], IN1[10], IN2);
  UB1BPPG_11_11 U11 (O[22], IN1[11], IN2);
  UB1BPPG_12_11 U12 (O[23], IN1[12], IN2);
  UB1BPPG_13_11 U13 (O[24], IN1[13], IN2);
  UB1BPPG_14_11 U14 (O[25], IN1[14], IN2);
  UB1BPPG_15_11 U15 (O[26], IN1[15], IN2);
endmodule

module UBVPPG_15_0_12 (O, IN1, IN2);
  output [27:12] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_12 U0 (O[12], IN1[0], IN2);
  UB1BPPG_1_12 U1 (O[13], IN1[1], IN2);
  UB1BPPG_2_12 U2 (O[14], IN1[2], IN2);
  UB1BPPG_3_12 U3 (O[15], IN1[3], IN2);
  UB1BPPG_4_12 U4 (O[16], IN1[4], IN2);
  UB1BPPG_5_12 U5 (O[17], IN1[5], IN2);
  UB1BPPG_6_12 U6 (O[18], IN1[6], IN2);
  UB1BPPG_7_12 U7 (O[19], IN1[7], IN2);
  UB1BPPG_8_12 U8 (O[20], IN1[8], IN2);
  UB1BPPG_9_12 U9 (O[21], IN1[9], IN2);
  UB1BPPG_10_12 U10 (O[22], IN1[10], IN2);
  UB1BPPG_11_12 U11 (O[23], IN1[11], IN2);
  UB1BPPG_12_12 U12 (O[24], IN1[12], IN2);
  UB1BPPG_13_12 U13 (O[25], IN1[13], IN2);
  UB1BPPG_14_12 U14 (O[26], IN1[14], IN2);
  UB1BPPG_15_12 U15 (O[27], IN1[15], IN2);
endmodule

module UBVPPG_15_0_13 (O, IN1, IN2);
  output [28:13] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_13 U0 (O[13], IN1[0], IN2);
  UB1BPPG_1_13 U1 (O[14], IN1[1], IN2);
  UB1BPPG_2_13 U2 (O[15], IN1[2], IN2);
  UB1BPPG_3_13 U3 (O[16], IN1[3], IN2);
  UB1BPPG_4_13 U4 (O[17], IN1[4], IN2);
  UB1BPPG_5_13 U5 (O[18], IN1[5], IN2);
  UB1BPPG_6_13 U6 (O[19], IN1[6], IN2);
  UB1BPPG_7_13 U7 (O[20], IN1[7], IN2);
  UB1BPPG_8_13 U8 (O[21], IN1[8], IN2);
  UB1BPPG_9_13 U9 (O[22], IN1[9], IN2);
  UB1BPPG_10_13 U10 (O[23], IN1[10], IN2);
  UB1BPPG_11_13 U11 (O[24], IN1[11], IN2);
  UB1BPPG_12_13 U12 (O[25], IN1[12], IN2);
  UB1BPPG_13_13 U13 (O[26], IN1[13], IN2);
  UB1BPPG_14_13 U14 (O[27], IN1[14], IN2);
  UB1BPPG_15_13 U15 (O[28], IN1[15], IN2);
endmodule

module UBVPPG_15_0_14 (O, IN1, IN2);
  output [29:14] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_14 U0 (O[14], IN1[0], IN2);
  UB1BPPG_1_14 U1 (O[15], IN1[1], IN2);
  UB1BPPG_2_14 U2 (O[16], IN1[2], IN2);
  UB1BPPG_3_14 U3 (O[17], IN1[3], IN2);
  UB1BPPG_4_14 U4 (O[18], IN1[4], IN2);
  UB1BPPG_5_14 U5 (O[19], IN1[5], IN2);
  UB1BPPG_6_14 U6 (O[20], IN1[6], IN2);
  UB1BPPG_7_14 U7 (O[21], IN1[7], IN2);
  UB1BPPG_8_14 U8 (O[22], IN1[8], IN2);
  UB1BPPG_9_14 U9 (O[23], IN1[9], IN2);
  UB1BPPG_10_14 U10 (O[24], IN1[10], IN2);
  UB1BPPG_11_14 U11 (O[25], IN1[11], IN2);
  UB1BPPG_12_14 U12 (O[26], IN1[12], IN2);
  UB1BPPG_13_14 U13 (O[27], IN1[13], IN2);
  UB1BPPG_14_14 U14 (O[28], IN1[14], IN2);
  UB1BPPG_15_14 U15 (O[29], IN1[15], IN2);
endmodule

module UBVPPG_15_0_15 (O, IN1, IN2);
  output [30:15] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_15 U0 (O[15], IN1[0], IN2);
  UB1BPPG_1_15 U1 (O[16], IN1[1], IN2);
  UB1BPPG_2_15 U2 (O[17], IN1[2], IN2);
  UB1BPPG_3_15 U3 (O[18], IN1[3], IN2);
  UB1BPPG_4_15 U4 (O[19], IN1[4], IN2);
  UB1BPPG_5_15 U5 (O[20], IN1[5], IN2);
  UB1BPPG_6_15 U6 (O[21], IN1[6], IN2);
  UB1BPPG_7_15 U7 (O[22], IN1[7], IN2);
  UB1BPPG_8_15 U8 (O[23], IN1[8], IN2);
  UB1BPPG_9_15 U9 (O[24], IN1[9], IN2);
  UB1BPPG_10_15 U10 (O[25], IN1[10], IN2);
  UB1BPPG_11_15 U11 (O[26], IN1[11], IN2);
  UB1BPPG_12_15 U12 (O[27], IN1[12], IN2);
  UB1BPPG_13_15 U13 (O[28], IN1[13], IN2);
  UB1BPPG_14_15 U14 (O[29], IN1[14], IN2);
  UB1BPPG_15_15 U15 (O[30], IN1[15], IN2);
endmodule

module UBVPPG_15_0_2 (O, IN1, IN2);
  output [17:2] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_2 U0 (O[2], IN1[0], IN2);
  UB1BPPG_1_2 U1 (O[3], IN1[1], IN2);
  UB1BPPG_2_2 U2 (O[4], IN1[2], IN2);
  UB1BPPG_3_2 U3 (O[5], IN1[3], IN2);
  UB1BPPG_4_2 U4 (O[6], IN1[4], IN2);
  UB1BPPG_5_2 U5 (O[7], IN1[5], IN2);
  UB1BPPG_6_2 U6 (O[8], IN1[6], IN2);
  UB1BPPG_7_2 U7 (O[9], IN1[7], IN2);
  UB1BPPG_8_2 U8 (O[10], IN1[8], IN2);
  UB1BPPG_9_2 U9 (O[11], IN1[9], IN2);
  UB1BPPG_10_2 U10 (O[12], IN1[10], IN2);
  UB1BPPG_11_2 U11 (O[13], IN1[11], IN2);
  UB1BPPG_12_2 U12 (O[14], IN1[12], IN2);
  UB1BPPG_13_2 U13 (O[15], IN1[13], IN2);
  UB1BPPG_14_2 U14 (O[16], IN1[14], IN2);
  UB1BPPG_15_2 U15 (O[17], IN1[15], IN2);
endmodule

module UBVPPG_15_0_3 (O, IN1, IN2);
  output [18:3] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_3 U0 (O[3], IN1[0], IN2);
  UB1BPPG_1_3 U1 (O[4], IN1[1], IN2);
  UB1BPPG_2_3 U2 (O[5], IN1[2], IN2);
  UB1BPPG_3_3 U3 (O[6], IN1[3], IN2);
  UB1BPPG_4_3 U4 (O[7], IN1[4], IN2);
  UB1BPPG_5_3 U5 (O[8], IN1[5], IN2);
  UB1BPPG_6_3 U6 (O[9], IN1[6], IN2);
  UB1BPPG_7_3 U7 (O[10], IN1[7], IN2);
  UB1BPPG_8_3 U8 (O[11], IN1[8], IN2);
  UB1BPPG_9_3 U9 (O[12], IN1[9], IN2);
  UB1BPPG_10_3 U10 (O[13], IN1[10], IN2);
  UB1BPPG_11_3 U11 (O[14], IN1[11], IN2);
  UB1BPPG_12_3 U12 (O[15], IN1[12], IN2);
  UB1BPPG_13_3 U13 (O[16], IN1[13], IN2);
  UB1BPPG_14_3 U14 (O[17], IN1[14], IN2);
  UB1BPPG_15_3 U15 (O[18], IN1[15], IN2);
endmodule

module UBVPPG_15_0_4 (O, IN1, IN2);
  output [19:4] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_4 U0 (O[4], IN1[0], IN2);
  UB1BPPG_1_4 U1 (O[5], IN1[1], IN2);
  UB1BPPG_2_4 U2 (O[6], IN1[2], IN2);
  UB1BPPG_3_4 U3 (O[7], IN1[3], IN2);
  UB1BPPG_4_4 U4 (O[8], IN1[4], IN2);
  UB1BPPG_5_4 U5 (O[9], IN1[5], IN2);
  UB1BPPG_6_4 U6 (O[10], IN1[6], IN2);
  UB1BPPG_7_4 U7 (O[11], IN1[7], IN2);
  UB1BPPG_8_4 U8 (O[12], IN1[8], IN2);
  UB1BPPG_9_4 U9 (O[13], IN1[9], IN2);
  UB1BPPG_10_4 U10 (O[14], IN1[10], IN2);
  UB1BPPG_11_4 U11 (O[15], IN1[11], IN2);
  UB1BPPG_12_4 U12 (O[16], IN1[12], IN2);
  UB1BPPG_13_4 U13 (O[17], IN1[13], IN2);
  UB1BPPG_14_4 U14 (O[18], IN1[14], IN2);
  UB1BPPG_15_4 U15 (O[19], IN1[15], IN2);
endmodule

module UBVPPG_15_0_5 (O, IN1, IN2);
  output [20:5] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_5 U0 (O[5], IN1[0], IN2);
  UB1BPPG_1_5 U1 (O[6], IN1[1], IN2);
  UB1BPPG_2_5 U2 (O[7], IN1[2], IN2);
  UB1BPPG_3_5 U3 (O[8], IN1[3], IN2);
  UB1BPPG_4_5 U4 (O[9], IN1[4], IN2);
  UB1BPPG_5_5 U5 (O[10], IN1[5], IN2);
  UB1BPPG_6_5 U6 (O[11], IN1[6], IN2);
  UB1BPPG_7_5 U7 (O[12], IN1[7], IN2);
  UB1BPPG_8_5 U8 (O[13], IN1[8], IN2);
  UB1BPPG_9_5 U9 (O[14], IN1[9], IN2);
  UB1BPPG_10_5 U10 (O[15], IN1[10], IN2);
  UB1BPPG_11_5 U11 (O[16], IN1[11], IN2);
  UB1BPPG_12_5 U12 (O[17], IN1[12], IN2);
  UB1BPPG_13_5 U13 (O[18], IN1[13], IN2);
  UB1BPPG_14_5 U14 (O[19], IN1[14], IN2);
  UB1BPPG_15_5 U15 (O[20], IN1[15], IN2);
endmodule

module UBVPPG_15_0_6 (O, IN1, IN2);
  output [21:6] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_6 U0 (O[6], IN1[0], IN2);
  UB1BPPG_1_6 U1 (O[7], IN1[1], IN2);
  UB1BPPG_2_6 U2 (O[8], IN1[2], IN2);
  UB1BPPG_3_6 U3 (O[9], IN1[3], IN2);
  UB1BPPG_4_6 U4 (O[10], IN1[4], IN2);
  UB1BPPG_5_6 U5 (O[11], IN1[5], IN2);
  UB1BPPG_6_6 U6 (O[12], IN1[6], IN2);
  UB1BPPG_7_6 U7 (O[13], IN1[7], IN2);
  UB1BPPG_8_6 U8 (O[14], IN1[8], IN2);
  UB1BPPG_9_6 U9 (O[15], IN1[9], IN2);
  UB1BPPG_10_6 U10 (O[16], IN1[10], IN2);
  UB1BPPG_11_6 U11 (O[17], IN1[11], IN2);
  UB1BPPG_12_6 U12 (O[18], IN1[12], IN2);
  UB1BPPG_13_6 U13 (O[19], IN1[13], IN2);
  UB1BPPG_14_6 U14 (O[20], IN1[14], IN2);
  UB1BPPG_15_6 U15 (O[21], IN1[15], IN2);
endmodule

module UBVPPG_15_0_7 (O, IN1, IN2);
  output [22:7] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_7 U0 (O[7], IN1[0], IN2);
  UB1BPPG_1_7 U1 (O[8], IN1[1], IN2);
  UB1BPPG_2_7 U2 (O[9], IN1[2], IN2);
  UB1BPPG_3_7 U3 (O[10], IN1[3], IN2);
  UB1BPPG_4_7 U4 (O[11], IN1[4], IN2);
  UB1BPPG_5_7 U5 (O[12], IN1[5], IN2);
  UB1BPPG_6_7 U6 (O[13], IN1[6], IN2);
  UB1BPPG_7_7 U7 (O[14], IN1[7], IN2);
  UB1BPPG_8_7 U8 (O[15], IN1[8], IN2);
  UB1BPPG_9_7 U9 (O[16], IN1[9], IN2);
  UB1BPPG_10_7 U10 (O[17], IN1[10], IN2);
  UB1BPPG_11_7 U11 (O[18], IN1[11], IN2);
  UB1BPPG_12_7 U12 (O[19], IN1[12], IN2);
  UB1BPPG_13_7 U13 (O[20], IN1[13], IN2);
  UB1BPPG_14_7 U14 (O[21], IN1[14], IN2);
  UB1BPPG_15_7 U15 (O[22], IN1[15], IN2);
endmodule

module UBVPPG_15_0_8 (O, IN1, IN2);
  output [23:8] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_8 U0 (O[8], IN1[0], IN2);
  UB1BPPG_1_8 U1 (O[9], IN1[1], IN2);
  UB1BPPG_2_8 U2 (O[10], IN1[2], IN2);
  UB1BPPG_3_8 U3 (O[11], IN1[3], IN2);
  UB1BPPG_4_8 U4 (O[12], IN1[4], IN2);
  UB1BPPG_5_8 U5 (O[13], IN1[5], IN2);
  UB1BPPG_6_8 U6 (O[14], IN1[6], IN2);
  UB1BPPG_7_8 U7 (O[15], IN1[7], IN2);
  UB1BPPG_8_8 U8 (O[16], IN1[8], IN2);
  UB1BPPG_9_8 U9 (O[17], IN1[9], IN2);
  UB1BPPG_10_8 U10 (O[18], IN1[10], IN2);
  UB1BPPG_11_8 U11 (O[19], IN1[11], IN2);
  UB1BPPG_12_8 U12 (O[20], IN1[12], IN2);
  UB1BPPG_13_8 U13 (O[21], IN1[13], IN2);
  UB1BPPG_14_8 U14 (O[22], IN1[14], IN2);
  UB1BPPG_15_8 U15 (O[23], IN1[15], IN2);
endmodule

module UBVPPG_15_0_9 (O, IN1, IN2);
  output [24:9] O;
  input [15:0] IN1;
  input IN2;
  UB1BPPG_0_9 U0 (O[9], IN1[0], IN2);
  UB1BPPG_1_9 U1 (O[10], IN1[1], IN2);
  UB1BPPG_2_9 U2 (O[11], IN1[2], IN2);
  UB1BPPG_3_9 U3 (O[12], IN1[3], IN2);
  UB1BPPG_4_9 U4 (O[13], IN1[4], IN2);
  UB1BPPG_5_9 U5 (O[14], IN1[5], IN2);
  UB1BPPG_6_9 U6 (O[15], IN1[6], IN2);
  UB1BPPG_7_9 U7 (O[16], IN1[7], IN2);
  UB1BPPG_8_9 U8 (O[17], IN1[8], IN2);
  UB1BPPG_9_9 U9 (O[18], IN1[9], IN2);
  UB1BPPG_10_9 U10 (O[19], IN1[10], IN2);
  UB1BPPG_11_9 U11 (O[20], IN1[11], IN2);
  UB1BPPG_12_9 U12 (O[21], IN1[12], IN2);
  UB1BPPG_13_9 U13 (O[22], IN1[13], IN2);
  UB1BPPG_14_9 U14 (O[23], IN1[14], IN2);
  UB1BPPG_15_9 U15 (O[24], IN1[15], IN2);
endmodule

